VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO regfile
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN regfile 0 0 ;
  SIZE 95.8 BY 1.55 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 95.8 1.75 ;
        RECT 95.485 1.045 95.55 1.75 ;
        RECT 94.73 1.045 94.795 1.75 ;
        RECT 94.385 1.045 94.45 1.75 ;
        RECT 93.83 1.045 93.895 1.75 ;
        RECT 93.455 1.045 93.52 1.75 ;
        RECT 92.7 1.045 92.765 1.75 ;
        RECT 92.355 1.045 92.42 1.75 ;
        RECT 91.8 1.045 91.865 1.75 ;
        RECT 90.5025 1.3475 91.0825 1.75 ;
        RECT 90.1925 1.045 90.2575 1.75 ;
        RECT 88.895 1.3475 89.475 1.75 ;
        RECT 88.585 1.045 88.65 1.75 ;
        RECT 88.215 1.045 88.28 1.75 ;
        RECT 85.9875 1.3475 87.225 1.75 ;
        RECT 85.6775 1.045 85.7425 1.75 ;
        RECT 85.3075 1.045 85.3725 1.75 ;
        RECT 83.08 1.3475 84.3175 1.75 ;
        RECT 82.77 1.045 82.835 1.75 ;
        RECT 82.4 1.045 82.465 1.75 ;
        RECT 80.1725 1.3475 81.41 1.75 ;
        RECT 79.8625 1.045 79.9275 1.75 ;
        RECT 79.4925 1.045 79.5575 1.75 ;
        RECT 77.265 1.3475 78.5025 1.75 ;
        RECT 76.955 1.045 77.02 1.75 ;
        RECT 76.585 1.045 76.65 1.75 ;
        RECT 74.3575 1.3475 75.595 1.75 ;
        RECT 74.0475 1.045 74.1125 1.75 ;
        RECT 73.6775 1.045 73.7425 1.75 ;
        RECT 71.45 1.3475 72.6875 1.75 ;
        RECT 71.14 1.045 71.205 1.75 ;
        RECT 70.77 1.045 70.835 1.75 ;
        RECT 68.5425 1.3475 69.78 1.75 ;
        RECT 68.2325 1.045 68.2975 1.75 ;
        RECT 67.8625 1.045 67.9275 1.75 ;
        RECT 65.635 1.3475 66.8725 1.75 ;
        RECT 65.325 1.045 65.39 1.75 ;
        RECT 64.955 1.045 65.02 1.75 ;
        RECT 62.7275 1.3475 63.965 1.75 ;
        RECT 62.4175 1.045 62.4825 1.75 ;
        RECT 62.0475 1.045 62.1125 1.75 ;
        RECT 59.82 1.3475 61.0575 1.75 ;
        RECT 59.51 1.045 59.575 1.75 ;
        RECT 59.14 1.045 59.205 1.75 ;
        RECT 56.9125 1.3475 58.15 1.75 ;
        RECT 56.6025 1.045 56.6675 1.75 ;
        RECT 56.2325 1.045 56.2975 1.75 ;
        RECT 54.005 1.3475 55.2425 1.75 ;
        RECT 53.695 1.045 53.76 1.75 ;
        RECT 53.325 1.045 53.39 1.75 ;
        RECT 51.0975 1.3475 52.335 1.75 ;
        RECT 50.7875 1.045 50.8525 1.75 ;
        RECT 50.4175 1.045 50.4825 1.75 ;
        RECT 48.19 1.3475 49.4275 1.75 ;
        RECT 47.88 1.045 47.945 1.75 ;
        RECT 47.51 1.045 47.575 1.75 ;
        RECT 45.2825 1.3475 46.52 1.75 ;
        RECT 44.9725 1.045 45.0375 1.75 ;
        RECT 44.6025 1.045 44.6675 1.75 ;
        RECT 42.375 1.3475 43.6125 1.75 ;
        RECT 42.065 1.045 42.13 1.75 ;
        RECT 41.695 1.045 41.76 1.75 ;
        RECT 39.4675 1.3475 40.705 1.75 ;
        RECT 39.1575 1.045 39.2225 1.75 ;
        RECT 38.7875 1.045 38.8525 1.75 ;
        RECT 36.56 1.3475 37.7975 1.75 ;
        RECT 36.25 1.045 36.315 1.75 ;
        RECT 35.88 1.045 35.945 1.75 ;
        RECT 33.6525 1.3475 34.89 1.75 ;
        RECT 33.3425 1.045 33.4075 1.75 ;
        RECT 32.9725 1.045 33.0375 1.75 ;
        RECT 30.745 1.3475 31.9825 1.75 ;
        RECT 30.435 1.045 30.5 1.75 ;
        RECT 30.065 1.045 30.13 1.75 ;
        RECT 27.8375 1.3475 29.075 1.75 ;
        RECT 27.5275 1.045 27.5925 1.75 ;
        RECT 27.1575 1.045 27.2225 1.75 ;
        RECT 24.93 1.3475 26.1675 1.75 ;
        RECT 24.62 1.045 24.685 1.75 ;
        RECT 24.25 1.045 24.315 1.75 ;
        RECT 22.0225 1.3475 23.26 1.75 ;
        RECT 21.7125 1.045 21.7775 1.75 ;
        RECT 21.3425 1.045 21.4075 1.75 ;
        RECT 19.115 1.3475 20.3525 1.75 ;
        RECT 18.805 1.045 18.87 1.75 ;
        RECT 18.435 1.045 18.5 1.75 ;
        RECT 16.2075 1.3475 17.445 1.75 ;
        RECT 15.8975 1.045 15.9625 1.75 ;
        RECT 15.5275 1.045 15.5925 1.75 ;
        RECT 13.3 1.3475 14.5375 1.75 ;
        RECT 12.99 1.045 13.055 1.75 ;
        RECT 12.62 1.045 12.685 1.75 ;
        RECT 10.3925 1.3475 11.63 1.75 ;
        RECT 10.0825 1.045 10.1475 1.75 ;
        RECT 9.7125 1.045 9.7775 1.75 ;
        RECT 7.485 1.3475 8.7225 1.75 ;
        RECT 7.175 1.045 7.24 1.75 ;
        RECT 6.805 1.045 6.87 1.75 ;
        RECT 4.5775 1.3475 5.815 1.75 ;
        RECT 4.2675 1.045 4.3325 1.75 ;
        RECT 3.8975 1.045 3.9625 1.75 ;
        RECT 1.67 1.3475 2.9075 1.75 ;
        RECT 1.36 1.045 1.425 1.75 ;
        RECT 0.99 1.045 1.055 1.75 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.2 95.8 0.2 ;
        RECT 95.485 -0.2 95.55 0.4225 ;
        RECT 94.73 -0.2 94.795 0.4225 ;
        RECT 94.385 -0.2 94.45 0.4225 ;
        RECT 93.83 -0.2 93.895 0.4225 ;
        RECT 93.455 -0.2 93.52 0.4225 ;
        RECT 92.7 -0.2 92.765 0.4225 ;
        RECT 92.355 -0.2 92.42 0.4225 ;
        RECT 91.8 -0.2 91.865 0.4225 ;
        RECT 90.1775 0.7875 90.3125 0.8525 ;
        RECT 90.1925 -0.2 90.2575 0.8525 ;
        RECT 88.585 -0.2 88.65 0.4225 ;
        RECT 88.215 -0.2 88.28 0.4225 ;
        RECT 85.6775 -0.2 85.7425 0.4225 ;
        RECT 85.3075 -0.2 85.3725 0.4225 ;
        RECT 82.77 -0.2 82.835 0.4225 ;
        RECT 82.4 -0.2 82.465 0.4225 ;
        RECT 79.8625 -0.2 79.9275 0.4225 ;
        RECT 79.4925 -0.2 79.5575 0.4225 ;
        RECT 76.955 -0.2 77.02 0.4225 ;
        RECT 76.585 -0.2 76.65 0.4225 ;
        RECT 74.0475 -0.2 74.1125 0.4225 ;
        RECT 73.6775 -0.2 73.7425 0.4225 ;
        RECT 71.14 -0.2 71.205 0.4225 ;
        RECT 70.77 -0.2 70.835 0.4225 ;
        RECT 68.2325 -0.2 68.2975 0.4225 ;
        RECT 67.8625 -0.2 67.9275 0.4225 ;
        RECT 65.325 -0.2 65.39 0.4225 ;
        RECT 64.955 -0.2 65.02 0.4225 ;
        RECT 62.4175 -0.2 62.4825 0.4225 ;
        RECT 62.0475 -0.2 62.1125 0.4225 ;
        RECT 59.51 -0.2 59.575 0.4225 ;
        RECT 59.14 -0.2 59.205 0.4225 ;
        RECT 56.6025 -0.2 56.6675 0.4225 ;
        RECT 56.2325 -0.2 56.2975 0.4225 ;
        RECT 53.695 -0.2 53.76 0.4225 ;
        RECT 53.325 -0.2 53.39 0.4225 ;
        RECT 50.7875 -0.2 50.8525 0.4225 ;
        RECT 50.4175 -0.2 50.4825 0.4225 ;
        RECT 47.88 -0.2 47.945 0.4225 ;
        RECT 47.51 -0.2 47.575 0.4225 ;
        RECT 44.9725 -0.2 45.0375 0.4225 ;
        RECT 44.6025 -0.2 44.6675 0.4225 ;
        RECT 42.065 -0.2 42.13 0.4225 ;
        RECT 41.695 -0.2 41.76 0.4225 ;
        RECT 39.1575 -0.2 39.2225 0.4225 ;
        RECT 38.7875 -0.2 38.8525 0.4225 ;
        RECT 36.25 -0.2 36.315 0.4225 ;
        RECT 35.88 -0.2 35.945 0.4225 ;
        RECT 33.3425 -0.2 33.4075 0.4225 ;
        RECT 32.9725 -0.2 33.0375 0.4225 ;
        RECT 30.435 -0.2 30.5 0.4225 ;
        RECT 30.065 -0.2 30.13 0.4225 ;
        RECT 27.5275 -0.2 27.5925 0.4225 ;
        RECT 27.1575 -0.2 27.2225 0.4225 ;
        RECT 24.62 -0.2 24.685 0.4225 ;
        RECT 24.25 -0.2 24.315 0.4225 ;
        RECT 21.7125 -0.2 21.7775 0.4225 ;
        RECT 21.3425 -0.2 21.4075 0.4225 ;
        RECT 18.805 -0.2 18.87 0.4225 ;
        RECT 18.435 -0.2 18.5 0.4225 ;
        RECT 15.8975 -0.2 15.9625 0.4225 ;
        RECT 15.5275 -0.2 15.5925 0.4225 ;
        RECT 12.99 -0.2 13.055 0.4225 ;
        RECT 12.62 -0.2 12.685 0.4225 ;
        RECT 10.0825 -0.2 10.1475 0.4225 ;
        RECT 9.7125 -0.2 9.7775 0.4225 ;
        RECT 7.175 -0.2 7.24 0.4225 ;
        RECT 6.805 -0.2 6.87 0.4225 ;
        RECT 4.2675 -0.2 4.3325 0.4225 ;
        RECT 3.8975 -0.2 3.9625 0.4225 ;
        RECT 1.36 -0.2 1.425 0.4225 ;
        RECT 0.99 -0.2 1.055 0.4225 ;
    END
  END vss!
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 94.34 0.7075 94.41 0.8425 ;
        RECT 92.31 0.7075 92.38 0.8425 ;
      LAYER metal2 ;
        RECT 92.27 0.1175 94.445 0.1875 ;
        RECT 94.34 0.705 94.41 0.845 ;
        RECT 92.31 0.705 92.38 0.845 ;
      LAYER metal3 ;
        RECT 94.305 0.1175 94.445 0.1875 ;
        RECT 94.34 0.055 94.41 1.4925 ;
        RECT 92.27 0.1175 92.41 0.1875 ;
        RECT 92.31 0.055 92.38 1.4925 ;
      LAYER via1 ;
        RECT 92.3125 0.7425 92.3775 0.8075 ;
        RECT 94.3425 0.7425 94.4075 0.8075 ;
      LAYER via2 ;
        RECT 92.305 0.1175 92.375 0.1875 ;
        RECT 92.31 0.74 92.38 0.81 ;
        RECT 94.34 0.74 94.41 0.81 ;
        RECT 94.34 0.1175 94.41 0.1875 ;
    END
  END clk
  PIN rd_mux_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.12 0.6975 87.485 0.8375 ;
      LAYER metal4 ;
        RECT 87.345 0.6975 87.485 0.8375 ;
        RECT 84.4375 0.6975 84.5775 0.8375 ;
        RECT 81.53 0.6975 81.67 0.8375 ;
        RECT 78.6225 0.6975 78.7625 0.8375 ;
        RECT 75.715 0.6975 75.855 0.8375 ;
        RECT 72.8075 0.6975 72.9475 0.8375 ;
        RECT 69.9 0.6975 70.04 0.8375 ;
        RECT 66.9925 0.6975 67.1325 0.8375 ;
        RECT 64.085 0.6975 64.225 0.8375 ;
        RECT 61.1775 0.6975 61.3175 0.8375 ;
        RECT 58.27 0.6975 58.41 0.8375 ;
        RECT 55.3625 0.6975 55.5025 0.8375 ;
        RECT 52.455 0.6975 52.595 0.8375 ;
        RECT 49.5475 0.6975 49.6875 0.8375 ;
        RECT 46.64 0.6975 46.78 0.8375 ;
        RECT 43.7325 0.6975 43.8725 0.8375 ;
        RECT 40.825 0.6975 40.965 0.8375 ;
        RECT 37.9175 0.6975 38.0575 0.8375 ;
        RECT 35.01 0.6975 35.15 0.8375 ;
        RECT 32.1025 0.6975 32.2425 0.8375 ;
        RECT 29.195 0.6975 29.335 0.8375 ;
        RECT 26.2875 0.6975 26.4275 0.8375 ;
        RECT 23.38 0.6975 23.52 0.8375 ;
        RECT 20.4725 0.6975 20.6125 0.8375 ;
        RECT 17.565 0.6975 17.705 0.8375 ;
        RECT 14.6575 0.6975 14.7975 0.8375 ;
        RECT 11.75 0.6975 11.89 0.8375 ;
        RECT 8.8425 0.6975 8.9825 0.8375 ;
        RECT 5.935 0.6975 6.075 0.8375 ;
        RECT 3.0275 0.6975 3.1675 0.8375 ;
        RECT 0.12 0.6975 0.26 0.8375 ;
      LAYER metal1 ;
        RECT 87.38 0.2725 87.45 0.4075 ;
        RECT 87.3825 0.265 87.4475 0.415 ;
        RECT 87.38 1.095 87.45 1.23 ;
        RECT 87.3825 1.0425 87.4475 1.2825 ;
        RECT 84.4725 0.2725 84.5425 0.4075 ;
        RECT 84.475 0.265 84.54 0.415 ;
        RECT 84.4725 1.095 84.5425 1.23 ;
        RECT 84.475 1.0425 84.54 1.2825 ;
        RECT 81.565 0.2725 81.635 0.4075 ;
        RECT 81.5675 0.265 81.6325 0.415 ;
        RECT 81.565 1.095 81.635 1.23 ;
        RECT 81.5675 1.0425 81.6325 1.2825 ;
        RECT 78.6575 0.2725 78.7275 0.4075 ;
        RECT 78.66 0.265 78.725 0.415 ;
        RECT 78.6575 1.095 78.7275 1.23 ;
        RECT 78.66 1.0425 78.725 1.2825 ;
        RECT 75.75 0.2725 75.82 0.4075 ;
        RECT 75.7525 0.265 75.8175 0.415 ;
        RECT 75.75 1.095 75.82 1.23 ;
        RECT 75.7525 1.0425 75.8175 1.2825 ;
        RECT 72.8425 0.2725 72.9125 0.4075 ;
        RECT 72.845 0.265 72.91 0.415 ;
        RECT 72.8425 1.095 72.9125 1.23 ;
        RECT 72.845 1.0425 72.91 1.2825 ;
        RECT 69.935 0.2725 70.005 0.4075 ;
        RECT 69.9375 0.265 70.0025 0.415 ;
        RECT 69.935 1.095 70.005 1.23 ;
        RECT 69.9375 1.0425 70.0025 1.2825 ;
        RECT 67.0275 0.2725 67.0975 0.4075 ;
        RECT 67.03 0.265 67.095 0.415 ;
        RECT 67.0275 1.095 67.0975 1.23 ;
        RECT 67.03 1.0425 67.095 1.2825 ;
        RECT 64.12 0.2725 64.19 0.4075 ;
        RECT 64.1225 0.265 64.1875 0.415 ;
        RECT 64.12 1.095 64.19 1.23 ;
        RECT 64.1225 1.0425 64.1875 1.2825 ;
        RECT 61.2125 0.2725 61.2825 0.4075 ;
        RECT 61.215 0.265 61.28 0.415 ;
        RECT 61.2125 1.095 61.2825 1.23 ;
        RECT 61.215 1.0425 61.28 1.2825 ;
        RECT 58.305 0.2725 58.375 0.4075 ;
        RECT 58.3075 0.265 58.3725 0.415 ;
        RECT 58.305 1.095 58.375 1.23 ;
        RECT 58.3075 1.0425 58.3725 1.2825 ;
        RECT 55.3975 0.2725 55.4675 0.4075 ;
        RECT 55.4 0.265 55.465 0.415 ;
        RECT 55.3975 1.095 55.4675 1.23 ;
        RECT 55.4 1.0425 55.465 1.2825 ;
        RECT 52.49 0.2725 52.56 0.4075 ;
        RECT 52.4925 0.265 52.5575 0.415 ;
        RECT 52.49 1.095 52.56 1.23 ;
        RECT 52.4925 1.0425 52.5575 1.2825 ;
        RECT 49.5825 0.2725 49.6525 0.4075 ;
        RECT 49.585 0.265 49.65 0.415 ;
        RECT 49.5825 1.095 49.6525 1.23 ;
        RECT 49.585 1.0425 49.65 1.2825 ;
        RECT 46.675 0.2725 46.745 0.4075 ;
        RECT 46.6775 0.265 46.7425 0.415 ;
        RECT 46.675 1.095 46.745 1.23 ;
        RECT 46.6775 1.0425 46.7425 1.2825 ;
        RECT 43.7675 0.2725 43.8375 0.4075 ;
        RECT 43.77 0.265 43.835 0.415 ;
        RECT 43.7675 1.095 43.8375 1.23 ;
        RECT 43.77 1.0425 43.835 1.2825 ;
        RECT 40.86 0.2725 40.93 0.4075 ;
        RECT 40.8625 0.265 40.9275 0.415 ;
        RECT 40.86 1.095 40.93 1.23 ;
        RECT 40.8625 1.0425 40.9275 1.2825 ;
        RECT 37.9525 0.2725 38.0225 0.4075 ;
        RECT 37.955 0.265 38.02 0.415 ;
        RECT 37.9525 1.095 38.0225 1.23 ;
        RECT 37.955 1.0425 38.02 1.2825 ;
        RECT 35.045 0.2725 35.115 0.4075 ;
        RECT 35.0475 0.265 35.1125 0.415 ;
        RECT 35.045 1.095 35.115 1.23 ;
        RECT 35.0475 1.0425 35.1125 1.2825 ;
        RECT 32.1375 0.2725 32.2075 0.4075 ;
        RECT 32.14 0.265 32.205 0.415 ;
        RECT 32.1375 1.095 32.2075 1.23 ;
        RECT 32.14 1.0425 32.205 1.2825 ;
        RECT 29.23 0.2725 29.3 0.4075 ;
        RECT 29.2325 0.265 29.2975 0.415 ;
        RECT 29.23 1.095 29.3 1.23 ;
        RECT 29.2325 1.0425 29.2975 1.2825 ;
        RECT 26.3225 0.2725 26.3925 0.4075 ;
        RECT 26.325 0.265 26.39 0.415 ;
        RECT 26.3225 1.095 26.3925 1.23 ;
        RECT 26.325 1.0425 26.39 1.2825 ;
        RECT 23.415 0.2725 23.485 0.4075 ;
        RECT 23.4175 0.265 23.4825 0.415 ;
        RECT 23.415 1.095 23.485 1.23 ;
        RECT 23.4175 1.0425 23.4825 1.2825 ;
        RECT 20.5075 0.2725 20.5775 0.4075 ;
        RECT 20.51 0.265 20.575 0.415 ;
        RECT 20.5075 1.095 20.5775 1.23 ;
        RECT 20.51 1.0425 20.575 1.2825 ;
        RECT 17.6 0.2725 17.67 0.4075 ;
        RECT 17.6025 0.265 17.6675 0.415 ;
        RECT 17.6 1.095 17.67 1.23 ;
        RECT 17.6025 1.0425 17.6675 1.2825 ;
        RECT 14.6925 0.2725 14.7625 0.4075 ;
        RECT 14.695 0.265 14.76 0.415 ;
        RECT 14.6925 1.095 14.7625 1.23 ;
        RECT 14.695 1.0425 14.76 1.2825 ;
        RECT 11.785 0.2725 11.855 0.4075 ;
        RECT 11.7875 0.265 11.8525 0.415 ;
        RECT 11.785 1.095 11.855 1.23 ;
        RECT 11.7875 1.0425 11.8525 1.2825 ;
        RECT 8.8775 0.2725 8.9475 0.4075 ;
        RECT 8.88 0.265 8.945 0.415 ;
        RECT 8.8775 1.095 8.9475 1.23 ;
        RECT 8.88 1.0425 8.945 1.2825 ;
        RECT 5.97 0.2725 6.04 0.4075 ;
        RECT 5.9725 0.265 6.0375 0.415 ;
        RECT 5.97 1.095 6.04 1.23 ;
        RECT 5.9725 1.0425 6.0375 1.2825 ;
        RECT 3.0625 0.2725 3.1325 0.4075 ;
        RECT 3.065 0.265 3.13 0.415 ;
        RECT 3.0625 1.095 3.1325 1.23 ;
        RECT 3.065 1.0425 3.13 1.2825 ;
        RECT 0.155 0.2725 0.225 0.4075 ;
        RECT 0.1575 0.265 0.2225 0.415 ;
        RECT 0.155 1.095 0.225 1.23 ;
        RECT 0.1575 1.0425 0.2225 1.2825 ;
      LAYER metal2 ;
        RECT 87.38 0.27 87.45 0.41 ;
        RECT 87.38 1.0925 87.45 1.2325 ;
        RECT 84.4725 0.27 84.5425 0.41 ;
        RECT 84.4725 1.0925 84.5425 1.2325 ;
        RECT 81.565 0.27 81.635 0.41 ;
        RECT 81.565 1.0925 81.635 1.2325 ;
        RECT 78.6575 0.27 78.7275 0.41 ;
        RECT 78.6575 1.0925 78.7275 1.2325 ;
        RECT 75.75 0.27 75.82 0.41 ;
        RECT 75.75 1.0925 75.82 1.2325 ;
        RECT 72.8425 0.27 72.9125 0.41 ;
        RECT 72.8425 1.0925 72.9125 1.2325 ;
        RECT 69.935 0.27 70.005 0.41 ;
        RECT 69.935 1.0925 70.005 1.2325 ;
        RECT 67.0275 0.27 67.0975 0.41 ;
        RECT 67.0275 1.0925 67.0975 1.2325 ;
        RECT 64.12 0.27 64.19 0.41 ;
        RECT 64.12 1.0925 64.19 1.2325 ;
        RECT 61.2125 0.27 61.2825 0.41 ;
        RECT 61.2125 1.0925 61.2825 1.2325 ;
        RECT 58.305 0.27 58.375 0.41 ;
        RECT 58.305 1.0925 58.375 1.2325 ;
        RECT 55.3975 0.27 55.4675 0.41 ;
        RECT 55.3975 1.0925 55.4675 1.2325 ;
        RECT 52.49 0.27 52.56 0.41 ;
        RECT 52.49 1.0925 52.56 1.2325 ;
        RECT 49.5825 0.27 49.6525 0.41 ;
        RECT 49.5825 1.0925 49.6525 1.2325 ;
        RECT 46.675 0.27 46.745 0.41 ;
        RECT 46.675 1.0925 46.745 1.2325 ;
        RECT 43.7675 0.27 43.8375 0.41 ;
        RECT 43.7675 1.0925 43.8375 1.2325 ;
        RECT 40.86 0.27 40.93 0.41 ;
        RECT 40.86 1.0925 40.93 1.2325 ;
        RECT 37.9525 0.27 38.0225 0.41 ;
        RECT 37.9525 1.0925 38.0225 1.2325 ;
        RECT 35.045 0.27 35.115 0.41 ;
        RECT 35.045 1.0925 35.115 1.2325 ;
        RECT 32.1375 0.27 32.2075 0.41 ;
        RECT 32.1375 1.0925 32.2075 1.2325 ;
        RECT 29.23 0.27 29.3 0.41 ;
        RECT 29.23 1.0925 29.3 1.2325 ;
        RECT 26.3225 0.27 26.3925 0.41 ;
        RECT 26.3225 1.0925 26.3925 1.2325 ;
        RECT 23.415 0.27 23.485 0.41 ;
        RECT 23.415 1.0925 23.485 1.2325 ;
        RECT 20.5075 0.27 20.5775 0.41 ;
        RECT 20.5075 1.0925 20.5775 1.2325 ;
        RECT 17.6 0.27 17.67 0.41 ;
        RECT 17.6 1.0925 17.67 1.2325 ;
        RECT 14.6925 0.27 14.7625 0.41 ;
        RECT 14.6925 1.0925 14.7625 1.2325 ;
        RECT 11.785 0.27 11.855 0.41 ;
        RECT 11.785 1.0925 11.855 1.2325 ;
        RECT 8.8775 0.27 8.9475 0.41 ;
        RECT 8.8775 1.0925 8.9475 1.2325 ;
        RECT 5.97 0.27 6.04 0.41 ;
        RECT 5.97 1.0925 6.04 1.2325 ;
        RECT 3.0625 0.27 3.1325 0.41 ;
        RECT 3.0625 1.0925 3.1325 1.2325 ;
        RECT 0.155 0.27 0.225 0.41 ;
        RECT 0.155 1.0925 0.225 1.2325 ;
      LAYER metal3 ;
        RECT 87.38 0.055 87.45 1.4925 ;
        RECT 84.4725 0.055 84.5425 1.4925 ;
        RECT 81.565 0.055 81.635 1.4925 ;
        RECT 78.6575 0.055 78.7275 1.4925 ;
        RECT 75.75 0.055 75.82 1.4925 ;
        RECT 72.8425 0.055 72.9125 1.4925 ;
        RECT 69.935 0.055 70.005 1.4925 ;
        RECT 67.0275 0.055 67.0975 1.4925 ;
        RECT 64.12 0.055 64.19 1.4925 ;
        RECT 61.2125 0.055 61.2825 1.4925 ;
        RECT 58.305 0.055 58.375 1.4925 ;
        RECT 55.3975 0.055 55.4675 1.4925 ;
        RECT 52.49 0.055 52.56 1.4925 ;
        RECT 49.5825 0.055 49.6525 1.4925 ;
        RECT 46.675 0.055 46.745 1.4925 ;
        RECT 43.7675 0.055 43.8375 1.4925 ;
        RECT 40.86 0.055 40.93 1.4925 ;
        RECT 37.9525 0.055 38.0225 1.4925 ;
        RECT 35.045 0.055 35.115 1.4925 ;
        RECT 32.1375 0.055 32.2075 1.4925 ;
        RECT 29.23 0.055 29.3 1.4925 ;
        RECT 26.3225 0.055 26.3925 1.4925 ;
        RECT 23.415 0.055 23.485 1.4925 ;
        RECT 20.5075 0.055 20.5775 1.4925 ;
        RECT 17.6 0.055 17.67 1.4925 ;
        RECT 14.6925 0.055 14.7625 1.4925 ;
        RECT 11.785 0.055 11.855 1.4925 ;
        RECT 8.8775 0.055 8.9475 1.4925 ;
        RECT 5.97 0.055 6.04 1.4925 ;
        RECT 3.0625 0.055 3.1325 1.4925 ;
        RECT 0.155 0.055 0.225 1.49 ;
      LAYER via4 ;
        RECT 0.12 0.6975 0.26 0.8375 ;
        RECT 3.0275 0.6975 3.1675 0.8375 ;
        RECT 5.935 0.6975 6.075 0.8375 ;
        RECT 8.8425 0.6975 8.9825 0.8375 ;
        RECT 11.75 0.6975 11.89 0.8375 ;
        RECT 14.6575 0.6975 14.7975 0.8375 ;
        RECT 17.565 0.6975 17.705 0.8375 ;
        RECT 20.4725 0.6975 20.6125 0.8375 ;
        RECT 23.38 0.6975 23.52 0.8375 ;
        RECT 26.2875 0.6975 26.4275 0.8375 ;
        RECT 29.195 0.6975 29.335 0.8375 ;
        RECT 32.1025 0.6975 32.2425 0.8375 ;
        RECT 35.01 0.6975 35.15 0.8375 ;
        RECT 37.9175 0.6975 38.0575 0.8375 ;
        RECT 40.825 0.6975 40.965 0.8375 ;
        RECT 43.7325 0.6975 43.8725 0.8375 ;
        RECT 46.64 0.6975 46.78 0.8375 ;
        RECT 49.5475 0.6975 49.6875 0.8375 ;
        RECT 52.455 0.6975 52.595 0.8375 ;
        RECT 55.3625 0.6975 55.5025 0.8375 ;
        RECT 58.27 0.6975 58.41 0.8375 ;
        RECT 61.1775 0.6975 61.3175 0.8375 ;
        RECT 64.085 0.6975 64.225 0.8375 ;
        RECT 66.9925 0.6975 67.1325 0.8375 ;
        RECT 69.9 0.6975 70.04 0.8375 ;
        RECT 72.8075 0.6975 72.9475 0.8375 ;
        RECT 75.715 0.6975 75.855 0.8375 ;
        RECT 78.6225 0.6975 78.7625 0.8375 ;
        RECT 81.53 0.6975 81.67 0.8375 ;
        RECT 84.4375 0.6975 84.5775 0.8375 ;
        RECT 87.345 0.6975 87.485 0.8375 ;
      LAYER via3 ;
        RECT 0.155 0.7325 0.225 0.8025 ;
        RECT 3.0625 0.7325 3.1325 0.8025 ;
        RECT 5.97 0.7325 6.04 0.8025 ;
        RECT 8.8775 0.7325 8.9475 0.8025 ;
        RECT 11.785 0.7325 11.855 0.8025 ;
        RECT 14.6925 0.7325 14.7625 0.8025 ;
        RECT 17.6 0.7325 17.67 0.8025 ;
        RECT 20.5075 0.7325 20.5775 0.8025 ;
        RECT 23.415 0.7325 23.485 0.8025 ;
        RECT 26.3225 0.7325 26.3925 0.8025 ;
        RECT 29.23 0.7325 29.3 0.8025 ;
        RECT 32.1375 0.7325 32.2075 0.8025 ;
        RECT 35.045 0.7325 35.115 0.8025 ;
        RECT 37.9525 0.7325 38.0225 0.8025 ;
        RECT 40.86 0.7325 40.93 0.8025 ;
        RECT 43.7675 0.7325 43.8375 0.8025 ;
        RECT 46.675 0.7325 46.745 0.8025 ;
        RECT 49.5825 0.7325 49.6525 0.8025 ;
        RECT 52.49 0.7325 52.56 0.8025 ;
        RECT 55.3975 0.7325 55.4675 0.8025 ;
        RECT 58.305 0.7325 58.375 0.8025 ;
        RECT 61.2125 0.7325 61.2825 0.8025 ;
        RECT 64.12 0.7325 64.19 0.8025 ;
        RECT 67.0275 0.7325 67.0975 0.8025 ;
        RECT 69.935 0.7325 70.005 0.8025 ;
        RECT 72.8425 0.7325 72.9125 0.8025 ;
        RECT 75.75 0.7325 75.82 0.8025 ;
        RECT 78.6575 0.7325 78.7275 0.8025 ;
        RECT 81.565 0.7325 81.635 0.8025 ;
        RECT 84.4725 0.7325 84.5425 0.8025 ;
        RECT 87.38 0.7325 87.45 0.8025 ;
      LAYER via1 ;
        RECT 0.1575 1.13 0.2225 1.195 ;
        RECT 0.1575 0.3075 0.2225 0.3725 ;
        RECT 3.065 1.13 3.13 1.195 ;
        RECT 3.065 0.3075 3.13 0.3725 ;
        RECT 5.9725 1.13 6.0375 1.195 ;
        RECT 5.9725 0.3075 6.0375 0.3725 ;
        RECT 8.88 1.13 8.945 1.195 ;
        RECT 8.88 0.3075 8.945 0.3725 ;
        RECT 11.7875 1.13 11.8525 1.195 ;
        RECT 11.7875 0.3075 11.8525 0.3725 ;
        RECT 14.695 1.13 14.76 1.195 ;
        RECT 14.695 0.3075 14.76 0.3725 ;
        RECT 17.6025 1.13 17.6675 1.195 ;
        RECT 17.6025 0.3075 17.6675 0.3725 ;
        RECT 20.51 1.13 20.575 1.195 ;
        RECT 20.51 0.3075 20.575 0.3725 ;
        RECT 23.4175 1.13 23.4825 1.195 ;
        RECT 23.4175 0.3075 23.4825 0.3725 ;
        RECT 26.325 1.13 26.39 1.195 ;
        RECT 26.325 0.3075 26.39 0.3725 ;
        RECT 29.2325 1.13 29.2975 1.195 ;
        RECT 29.2325 0.3075 29.2975 0.3725 ;
        RECT 32.14 1.13 32.205 1.195 ;
        RECT 32.14 0.3075 32.205 0.3725 ;
        RECT 35.0475 1.13 35.1125 1.195 ;
        RECT 35.0475 0.3075 35.1125 0.3725 ;
        RECT 37.955 1.13 38.02 1.195 ;
        RECT 37.955 0.3075 38.02 0.3725 ;
        RECT 40.8625 1.13 40.9275 1.195 ;
        RECT 40.8625 0.3075 40.9275 0.3725 ;
        RECT 43.77 1.13 43.835 1.195 ;
        RECT 43.77 0.3075 43.835 0.3725 ;
        RECT 46.6775 1.13 46.7425 1.195 ;
        RECT 46.6775 0.3075 46.7425 0.3725 ;
        RECT 49.585 1.13 49.65 1.195 ;
        RECT 49.585 0.3075 49.65 0.3725 ;
        RECT 52.4925 1.13 52.5575 1.195 ;
        RECT 52.4925 0.3075 52.5575 0.3725 ;
        RECT 55.4 1.13 55.465 1.195 ;
        RECT 55.4 0.3075 55.465 0.3725 ;
        RECT 58.3075 1.13 58.3725 1.195 ;
        RECT 58.3075 0.3075 58.3725 0.3725 ;
        RECT 61.215 1.13 61.28 1.195 ;
        RECT 61.215 0.3075 61.28 0.3725 ;
        RECT 64.1225 1.13 64.1875 1.195 ;
        RECT 64.1225 0.3075 64.1875 0.3725 ;
        RECT 67.03 1.13 67.095 1.195 ;
        RECT 67.03 0.3075 67.095 0.3725 ;
        RECT 69.9375 1.13 70.0025 1.195 ;
        RECT 69.9375 0.3075 70.0025 0.3725 ;
        RECT 72.845 1.13 72.91 1.195 ;
        RECT 72.845 0.3075 72.91 0.3725 ;
        RECT 75.7525 1.13 75.8175 1.195 ;
        RECT 75.7525 0.3075 75.8175 0.3725 ;
        RECT 78.66 1.13 78.725 1.195 ;
        RECT 78.66 0.3075 78.725 0.3725 ;
        RECT 81.5675 1.13 81.6325 1.195 ;
        RECT 81.5675 0.3075 81.6325 0.3725 ;
        RECT 84.475 1.13 84.54 1.195 ;
        RECT 84.475 0.3075 84.54 0.3725 ;
        RECT 87.3825 1.13 87.4475 1.195 ;
        RECT 87.3825 0.3075 87.4475 0.3725 ;
      LAYER via2 ;
        RECT 0.155 1.1275 0.225 1.1975 ;
        RECT 0.155 0.305 0.225 0.375 ;
        RECT 3.0625 1.1275 3.1325 1.1975 ;
        RECT 3.0625 0.305 3.1325 0.375 ;
        RECT 5.97 1.1275 6.04 1.1975 ;
        RECT 5.97 0.305 6.04 0.375 ;
        RECT 8.8775 1.1275 8.9475 1.1975 ;
        RECT 8.8775 0.305 8.9475 0.375 ;
        RECT 11.785 1.1275 11.855 1.1975 ;
        RECT 11.785 0.305 11.855 0.375 ;
        RECT 14.6925 1.1275 14.7625 1.1975 ;
        RECT 14.6925 0.305 14.7625 0.375 ;
        RECT 17.6 1.1275 17.67 1.1975 ;
        RECT 17.6 0.305 17.67 0.375 ;
        RECT 20.5075 1.1275 20.5775 1.1975 ;
        RECT 20.5075 0.305 20.5775 0.375 ;
        RECT 23.415 1.1275 23.485 1.1975 ;
        RECT 23.415 0.305 23.485 0.375 ;
        RECT 26.3225 1.1275 26.3925 1.1975 ;
        RECT 26.3225 0.305 26.3925 0.375 ;
        RECT 29.23 1.1275 29.3 1.1975 ;
        RECT 29.23 0.305 29.3 0.375 ;
        RECT 32.1375 1.1275 32.2075 1.1975 ;
        RECT 32.1375 0.305 32.2075 0.375 ;
        RECT 35.045 1.1275 35.115 1.1975 ;
        RECT 35.045 0.305 35.115 0.375 ;
        RECT 37.9525 1.1275 38.0225 1.1975 ;
        RECT 37.9525 0.305 38.0225 0.375 ;
        RECT 40.86 1.1275 40.93 1.1975 ;
        RECT 40.86 0.305 40.93 0.375 ;
        RECT 43.7675 1.1275 43.8375 1.1975 ;
        RECT 43.7675 0.305 43.8375 0.375 ;
        RECT 46.675 1.1275 46.745 1.1975 ;
        RECT 46.675 0.305 46.745 0.375 ;
        RECT 49.5825 1.1275 49.6525 1.1975 ;
        RECT 49.5825 0.305 49.6525 0.375 ;
        RECT 52.49 1.1275 52.56 1.1975 ;
        RECT 52.49 0.305 52.56 0.375 ;
        RECT 55.3975 1.1275 55.4675 1.1975 ;
        RECT 55.3975 0.305 55.4675 0.375 ;
        RECT 58.305 1.1275 58.375 1.1975 ;
        RECT 58.305 0.305 58.375 0.375 ;
        RECT 61.2125 1.1275 61.2825 1.1975 ;
        RECT 61.2125 0.305 61.2825 0.375 ;
        RECT 64.12 1.1275 64.19 1.1975 ;
        RECT 64.12 0.305 64.19 0.375 ;
        RECT 67.0275 1.1275 67.0975 1.1975 ;
        RECT 67.0275 0.305 67.0975 0.375 ;
        RECT 69.935 1.1275 70.005 1.1975 ;
        RECT 69.935 0.305 70.005 0.375 ;
        RECT 72.8425 1.1275 72.9125 1.1975 ;
        RECT 72.8425 0.305 72.9125 0.375 ;
        RECT 75.75 1.1275 75.82 1.1975 ;
        RECT 75.75 0.305 75.82 0.375 ;
        RECT 78.6575 1.1275 78.7275 1.1975 ;
        RECT 78.6575 0.305 78.7275 0.375 ;
        RECT 81.565 1.1275 81.635 1.1975 ;
        RECT 81.565 0.305 81.635 0.375 ;
        RECT 84.4725 1.1275 84.5425 1.1975 ;
        RECT 84.4725 0.305 84.5425 0.375 ;
        RECT 87.38 1.1275 87.45 1.1975 ;
        RECT 87.38 0.305 87.45 0.375 ;
    END
  END rd_mux_out
  PIN rd_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 61.9175 0.45 61.9875 0.585 ;
        RECT 61.6425 0.9075 61.985 0.9725 ;
        RECT 61.92 0.4475 61.985 0.9725 ;
        RECT 61.2725 0.53 61.4075 0.595 ;
      LAYER metal2 ;
        RECT 61.9175 0.12 61.9875 0.5875 ;
        RECT 61.0575 0.12 61.9875 0.19 ;
        RECT 61.0575 0.5275 61.4075 0.5975 ;
        RECT 61.0575 0.12 61.1275 0.5975 ;
      LAYER metal3 ;
        RECT 61.9175 0.055 61.9875 1.4925 ;
      LAYER via1 ;
        RECT 61.3075 0.53 61.3725 0.595 ;
        RECT 61.92 0.485 61.985 0.55 ;
      LAYER via2 ;
        RECT 61.9175 0.4825 61.9875 0.5525 ;
    END
  END rd_sel[10]
  PIN rd_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 59.01 0.45 59.08 0.585 ;
        RECT 58.735 0.9075 59.0775 0.9725 ;
        RECT 59.0125 0.4475 59.0775 0.9725 ;
        RECT 58.365 0.53 58.5 0.595 ;
      LAYER metal2 ;
        RECT 59.01 0.12 59.08 0.5875 ;
        RECT 58.15 0.12 59.08 0.19 ;
        RECT 58.15 0.5275 58.5 0.5975 ;
        RECT 58.15 0.12 58.22 0.5975 ;
      LAYER metal3 ;
        RECT 59.01 0.055 59.08 1.4925 ;
      LAYER via1 ;
        RECT 58.4 0.53 58.465 0.595 ;
        RECT 59.0125 0.485 59.0775 0.55 ;
      LAYER via2 ;
        RECT 59.01 0.4825 59.08 0.5525 ;
    END
  END rd_sel[11]
  PIN rd_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 56.1025 0.45 56.1725 0.585 ;
        RECT 55.8275 0.9075 56.17 0.9725 ;
        RECT 56.105 0.4475 56.17 0.9725 ;
        RECT 55.4575 0.53 55.5925 0.595 ;
      LAYER metal2 ;
        RECT 56.1025 0.12 56.1725 0.5875 ;
        RECT 55.2425 0.12 56.1725 0.19 ;
        RECT 55.2425 0.5275 55.5925 0.5975 ;
        RECT 55.2425 0.12 55.3125 0.5975 ;
      LAYER metal3 ;
        RECT 56.1025 0.055 56.1725 1.4925 ;
      LAYER via1 ;
        RECT 55.4925 0.53 55.5575 0.595 ;
        RECT 56.105 0.485 56.17 0.55 ;
      LAYER via2 ;
        RECT 56.1025 0.4825 56.1725 0.5525 ;
    END
  END rd_sel[12]
  PIN rd_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 53.195 0.45 53.265 0.585 ;
        RECT 52.92 0.9075 53.2625 0.9725 ;
        RECT 53.1975 0.4475 53.2625 0.9725 ;
        RECT 52.55 0.53 52.685 0.595 ;
      LAYER metal2 ;
        RECT 53.195 0.12 53.265 0.5875 ;
        RECT 52.335 0.12 53.265 0.19 ;
        RECT 52.335 0.5275 52.685 0.5975 ;
        RECT 52.335 0.12 52.405 0.5975 ;
      LAYER metal3 ;
        RECT 53.195 0.055 53.265 1.4925 ;
      LAYER via1 ;
        RECT 52.585 0.53 52.65 0.595 ;
        RECT 53.1975 0.485 53.2625 0.55 ;
      LAYER via2 ;
        RECT 53.195 0.4825 53.265 0.5525 ;
    END
  END rd_sel[13]
  PIN rd_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 50.2875 0.45 50.3575 0.585 ;
        RECT 50.0125 0.9075 50.355 0.9725 ;
        RECT 50.29 0.4475 50.355 0.9725 ;
        RECT 49.6425 0.53 49.7775 0.595 ;
      LAYER metal2 ;
        RECT 50.2875 0.12 50.3575 0.5875 ;
        RECT 49.4275 0.12 50.3575 0.19 ;
        RECT 49.4275 0.5275 49.7775 0.5975 ;
        RECT 49.4275 0.12 49.4975 0.5975 ;
      LAYER metal3 ;
        RECT 50.2875 0.055 50.3575 1.4925 ;
      LAYER via1 ;
        RECT 49.6775 0.53 49.7425 0.595 ;
        RECT 50.29 0.485 50.355 0.55 ;
      LAYER via2 ;
        RECT 50.2875 0.4825 50.3575 0.5525 ;
    END
  END rd_sel[14]
  PIN rd_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 47.38 0.45 47.45 0.585 ;
        RECT 47.105 0.9075 47.4475 0.9725 ;
        RECT 47.3825 0.4475 47.4475 0.9725 ;
        RECT 46.735 0.53 46.87 0.595 ;
      LAYER metal2 ;
        RECT 47.38 0.12 47.45 0.5875 ;
        RECT 46.52 0.12 47.45 0.19 ;
        RECT 46.52 0.5275 46.87 0.5975 ;
        RECT 46.52 0.12 46.59 0.5975 ;
      LAYER metal3 ;
        RECT 47.38 0.055 47.45 1.4925 ;
      LAYER via1 ;
        RECT 46.77 0.53 46.835 0.595 ;
        RECT 47.3825 0.485 47.4475 0.55 ;
      LAYER via2 ;
        RECT 47.38 0.4825 47.45 0.5525 ;
    END
  END rd_sel[15]
  PIN rd_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 44.4725 0.45 44.5425 0.585 ;
        RECT 44.1975 0.9075 44.54 0.9725 ;
        RECT 44.475 0.4475 44.54 0.9725 ;
        RECT 43.8275 0.53 43.9625 0.595 ;
      LAYER metal2 ;
        RECT 44.4725 0.12 44.5425 0.5875 ;
        RECT 43.6125 0.12 44.5425 0.19 ;
        RECT 43.6125 0.5275 43.9625 0.5975 ;
        RECT 43.6125 0.12 43.6825 0.5975 ;
      LAYER metal3 ;
        RECT 44.4725 0.055 44.5425 1.4925 ;
      LAYER via1 ;
        RECT 43.8625 0.53 43.9275 0.595 ;
        RECT 44.475 0.485 44.54 0.55 ;
      LAYER via2 ;
        RECT 44.4725 0.4825 44.5425 0.5525 ;
    END
  END rd_sel[16]
  PIN rd_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 41.565 0.45 41.635 0.585 ;
        RECT 41.29 0.9075 41.6325 0.9725 ;
        RECT 41.5675 0.4475 41.6325 0.9725 ;
        RECT 40.92 0.53 41.055 0.595 ;
      LAYER metal2 ;
        RECT 41.565 0.12 41.635 0.5875 ;
        RECT 40.705 0.12 41.635 0.19 ;
        RECT 40.705 0.5275 41.055 0.5975 ;
        RECT 40.705 0.12 40.775 0.5975 ;
      LAYER metal3 ;
        RECT 41.565 0.055 41.635 1.4925 ;
      LAYER via1 ;
        RECT 40.955 0.53 41.02 0.595 ;
        RECT 41.5675 0.485 41.6325 0.55 ;
      LAYER via2 ;
        RECT 41.565 0.4825 41.635 0.5525 ;
    END
  END rd_sel[17]
  PIN rd_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 38.6575 0.45 38.7275 0.585 ;
        RECT 38.3825 0.9075 38.725 0.9725 ;
        RECT 38.66 0.4475 38.725 0.9725 ;
        RECT 38.0125 0.53 38.1475 0.595 ;
      LAYER metal2 ;
        RECT 38.6575 0.12 38.7275 0.5875 ;
        RECT 37.7975 0.12 38.7275 0.19 ;
        RECT 37.7975 0.5275 38.1475 0.5975 ;
        RECT 37.7975 0.12 37.8675 0.5975 ;
      LAYER metal3 ;
        RECT 38.6575 0.055 38.7275 1.4925 ;
      LAYER via1 ;
        RECT 38.0475 0.53 38.1125 0.595 ;
        RECT 38.66 0.485 38.725 0.55 ;
      LAYER via2 ;
        RECT 38.6575 0.4825 38.7275 0.5525 ;
    END
  END rd_sel[18]
  PIN rd_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 35.75 0.45 35.82 0.585 ;
        RECT 35.475 0.9075 35.8175 0.9725 ;
        RECT 35.7525 0.4475 35.8175 0.9725 ;
        RECT 35.105 0.53 35.24 0.595 ;
      LAYER metal2 ;
        RECT 35.75 0.12 35.82 0.5875 ;
        RECT 34.89 0.12 35.82 0.19 ;
        RECT 34.89 0.5275 35.24 0.5975 ;
        RECT 34.89 0.12 34.96 0.5975 ;
      LAYER metal3 ;
        RECT 35.75 0.055 35.82 1.4925 ;
      LAYER via1 ;
        RECT 35.14 0.53 35.205 0.595 ;
        RECT 35.7525 0.485 35.8175 0.55 ;
      LAYER via2 ;
        RECT 35.75 0.4825 35.82 0.5525 ;
    END
  END rd_sel[19]
  PIN rd_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 88.085 0.45 88.155 0.585 ;
        RECT 87.81 0.9075 88.1525 0.9725 ;
        RECT 88.0875 0.4475 88.1525 0.9725 ;
        RECT 87.44 0.53 87.575 0.595 ;
      LAYER metal2 ;
        RECT 88.085 0.12 88.155 0.5875 ;
        RECT 87.225 0.12 88.155 0.19 ;
        RECT 87.225 0.5275 87.575 0.5975 ;
        RECT 87.225 0.12 87.295 0.5975 ;
      LAYER metal3 ;
        RECT 88.085 0.055 88.155 1.4925 ;
      LAYER via1 ;
        RECT 87.475 0.53 87.54 0.595 ;
        RECT 88.0875 0.485 88.1525 0.55 ;
      LAYER via2 ;
        RECT 88.085 0.4825 88.155 0.5525 ;
    END
  END rd_sel[1]
  PIN rd_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 32.8425 0.45 32.9125 0.585 ;
        RECT 32.5675 0.9075 32.91 0.9725 ;
        RECT 32.845 0.4475 32.91 0.9725 ;
        RECT 32.1975 0.53 32.3325 0.595 ;
      LAYER metal2 ;
        RECT 32.8425 0.12 32.9125 0.5875 ;
        RECT 31.9825 0.12 32.9125 0.19 ;
        RECT 31.9825 0.5275 32.3325 0.5975 ;
        RECT 31.9825 0.12 32.0525 0.5975 ;
      LAYER metal3 ;
        RECT 32.8425 0.055 32.9125 1.4925 ;
      LAYER via1 ;
        RECT 32.2325 0.53 32.2975 0.595 ;
        RECT 32.845 0.485 32.91 0.55 ;
      LAYER via2 ;
        RECT 32.8425 0.4825 32.9125 0.5525 ;
    END
  END rd_sel[20]
  PIN rd_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 29.935 0.45 30.005 0.585 ;
        RECT 29.66 0.9075 30.0025 0.9725 ;
        RECT 29.9375 0.4475 30.0025 0.9725 ;
        RECT 29.29 0.53 29.425 0.595 ;
      LAYER metal2 ;
        RECT 29.935 0.12 30.005 0.5875 ;
        RECT 29.075 0.12 30.005 0.19 ;
        RECT 29.075 0.5275 29.425 0.5975 ;
        RECT 29.075 0.12 29.145 0.5975 ;
      LAYER metal3 ;
        RECT 29.935 0.055 30.005 1.4925 ;
      LAYER via1 ;
        RECT 29.325 0.53 29.39 0.595 ;
        RECT 29.9375 0.485 30.0025 0.55 ;
      LAYER via2 ;
        RECT 29.935 0.4825 30.005 0.5525 ;
    END
  END rd_sel[21]
  PIN rd_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 27.0275 0.45 27.0975 0.585 ;
        RECT 26.7525 0.9075 27.095 0.9725 ;
        RECT 27.03 0.4475 27.095 0.9725 ;
        RECT 26.3825 0.53 26.5175 0.595 ;
      LAYER metal2 ;
        RECT 27.0275 0.12 27.0975 0.5875 ;
        RECT 26.1675 0.12 27.0975 0.19 ;
        RECT 26.1675 0.5275 26.5175 0.5975 ;
        RECT 26.1675 0.12 26.2375 0.5975 ;
      LAYER metal3 ;
        RECT 27.0275 0.055 27.0975 1.4925 ;
      LAYER via1 ;
        RECT 26.4175 0.53 26.4825 0.595 ;
        RECT 27.03 0.485 27.095 0.55 ;
      LAYER via2 ;
        RECT 27.0275 0.4825 27.0975 0.5525 ;
    END
  END rd_sel[22]
  PIN rd_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 24.12 0.45 24.19 0.585 ;
        RECT 23.845 0.9075 24.1875 0.9725 ;
        RECT 24.1225 0.4475 24.1875 0.9725 ;
        RECT 23.475 0.53 23.61 0.595 ;
      LAYER metal2 ;
        RECT 24.12 0.12 24.19 0.5875 ;
        RECT 23.26 0.12 24.19 0.19 ;
        RECT 23.26 0.5275 23.61 0.5975 ;
        RECT 23.26 0.12 23.33 0.5975 ;
      LAYER metal3 ;
        RECT 24.12 0.055 24.19 1.4925 ;
      LAYER via1 ;
        RECT 23.51 0.53 23.575 0.595 ;
        RECT 24.1225 0.485 24.1875 0.55 ;
      LAYER via2 ;
        RECT 24.12 0.4825 24.19 0.5525 ;
    END
  END rd_sel[23]
  PIN rd_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 21.2125 0.45 21.2825 0.585 ;
        RECT 20.9375 0.9075 21.28 0.9725 ;
        RECT 21.215 0.4475 21.28 0.9725 ;
        RECT 20.5675 0.53 20.7025 0.595 ;
      LAYER metal2 ;
        RECT 21.2125 0.12 21.2825 0.5875 ;
        RECT 20.3525 0.12 21.2825 0.19 ;
        RECT 20.3525 0.5275 20.7025 0.5975 ;
        RECT 20.3525 0.12 20.4225 0.5975 ;
      LAYER metal3 ;
        RECT 21.2125 0.055 21.2825 1.4925 ;
      LAYER via1 ;
        RECT 20.6025 0.53 20.6675 0.595 ;
        RECT 21.215 0.485 21.28 0.55 ;
      LAYER via2 ;
        RECT 21.2125 0.4825 21.2825 0.5525 ;
    END
  END rd_sel[24]
  PIN rd_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 18.305 0.45 18.375 0.585 ;
        RECT 18.03 0.9075 18.3725 0.9725 ;
        RECT 18.3075 0.4475 18.3725 0.9725 ;
        RECT 17.66 0.53 17.795 0.595 ;
      LAYER metal2 ;
        RECT 18.305 0.12 18.375 0.5875 ;
        RECT 17.445 0.12 18.375 0.19 ;
        RECT 17.445 0.5275 17.795 0.5975 ;
        RECT 17.445 0.12 17.515 0.5975 ;
      LAYER metal3 ;
        RECT 18.305 0.055 18.375 1.4925 ;
      LAYER via1 ;
        RECT 17.695 0.53 17.76 0.595 ;
        RECT 18.3075 0.485 18.3725 0.55 ;
      LAYER via2 ;
        RECT 18.305 0.4825 18.375 0.5525 ;
    END
  END rd_sel[25]
  PIN rd_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.3975 0.45 15.4675 0.585 ;
        RECT 15.1225 0.9075 15.465 0.9725 ;
        RECT 15.4 0.4475 15.465 0.9725 ;
        RECT 14.7525 0.53 14.8875 0.595 ;
      LAYER metal2 ;
        RECT 15.3975 0.12 15.4675 0.5875 ;
        RECT 14.5375 0.12 15.4675 0.19 ;
        RECT 14.5375 0.5275 14.8875 0.5975 ;
        RECT 14.5375 0.12 14.6075 0.5975 ;
      LAYER metal3 ;
        RECT 15.3975 0.055 15.4675 1.4925 ;
      LAYER via1 ;
        RECT 14.7875 0.53 14.8525 0.595 ;
        RECT 15.4 0.485 15.465 0.55 ;
      LAYER via2 ;
        RECT 15.3975 0.4825 15.4675 0.5525 ;
    END
  END rd_sel[26]
  PIN rd_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.49 0.45 12.56 0.585 ;
        RECT 12.215 0.9075 12.5575 0.9725 ;
        RECT 12.4925 0.4475 12.5575 0.9725 ;
        RECT 11.845 0.53 11.98 0.595 ;
      LAYER metal2 ;
        RECT 12.49 0.12 12.56 0.5875 ;
        RECT 11.63 0.12 12.56 0.19 ;
        RECT 11.63 0.5275 11.98 0.5975 ;
        RECT 11.63 0.12 11.7 0.5975 ;
      LAYER metal3 ;
        RECT 12.49 0.055 12.56 1.4925 ;
      LAYER via1 ;
        RECT 11.88 0.53 11.945 0.595 ;
        RECT 12.4925 0.485 12.5575 0.55 ;
      LAYER via2 ;
        RECT 12.49 0.4825 12.56 0.5525 ;
    END
  END rd_sel[27]
  PIN rd_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.5825 0.45 9.6525 0.585 ;
        RECT 9.3075 0.9075 9.65 0.9725 ;
        RECT 9.585 0.4475 9.65 0.9725 ;
        RECT 8.9375 0.53 9.0725 0.595 ;
      LAYER metal2 ;
        RECT 9.5825 0.12 9.6525 0.5875 ;
        RECT 8.7225 0.12 9.6525 0.19 ;
        RECT 8.7225 0.5275 9.0725 0.5975 ;
        RECT 8.7225 0.12 8.7925 0.5975 ;
      LAYER metal3 ;
        RECT 9.5825 0.055 9.6525 1.4925 ;
      LAYER via1 ;
        RECT 8.9725 0.53 9.0375 0.595 ;
        RECT 9.585 0.485 9.65 0.55 ;
      LAYER via2 ;
        RECT 9.5825 0.4825 9.6525 0.5525 ;
    END
  END rd_sel[28]
  PIN rd_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.675 0.45 6.745 0.585 ;
        RECT 6.4 0.9075 6.7425 0.9725 ;
        RECT 6.6775 0.4475 6.7425 0.9725 ;
        RECT 6.03 0.53 6.165 0.595 ;
      LAYER metal2 ;
        RECT 6.675 0.12 6.745 0.5875 ;
        RECT 5.815 0.12 6.745 0.19 ;
        RECT 5.815 0.5275 6.165 0.5975 ;
        RECT 5.815 0.12 5.885 0.5975 ;
      LAYER metal3 ;
        RECT 6.675 0.055 6.745 1.4925 ;
      LAYER via1 ;
        RECT 6.065 0.53 6.13 0.595 ;
        RECT 6.6775 0.485 6.7425 0.55 ;
      LAYER via2 ;
        RECT 6.675 0.4825 6.745 0.5525 ;
    END
  END rd_sel[29]
  PIN rd_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 85.1775 0.45 85.2475 0.585 ;
        RECT 84.9025 0.9075 85.245 0.9725 ;
        RECT 85.18 0.4475 85.245 0.9725 ;
        RECT 84.5325 0.53 84.6675 0.595 ;
      LAYER metal2 ;
        RECT 85.1775 0.12 85.2475 0.5875 ;
        RECT 84.3175 0.12 85.2475 0.19 ;
        RECT 84.3175 0.5275 84.6675 0.5975 ;
        RECT 84.3175 0.12 84.3875 0.5975 ;
      LAYER metal3 ;
        RECT 85.1775 0.055 85.2475 1.4925 ;
      LAYER via1 ;
        RECT 84.5675 0.53 84.6325 0.595 ;
        RECT 85.18 0.485 85.245 0.55 ;
      LAYER via2 ;
        RECT 85.1775 0.4825 85.2475 0.5525 ;
    END
  END rd_sel[2]
  PIN rd_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.7675 0.45 3.8375 0.585 ;
        RECT 3.4925 0.9075 3.835 0.9725 ;
        RECT 3.77 0.4475 3.835 0.9725 ;
        RECT 3.1225 0.53 3.2575 0.595 ;
      LAYER metal2 ;
        RECT 3.7675 0.12 3.8375 0.5875 ;
        RECT 2.9075 0.12 3.8375 0.19 ;
        RECT 2.9075 0.5275 3.2575 0.5975 ;
        RECT 2.9075 0.12 2.9775 0.5975 ;
      LAYER metal3 ;
        RECT 3.7675 0.055 3.8375 1.4925 ;
      LAYER via1 ;
        RECT 3.1575 0.53 3.2225 0.595 ;
        RECT 3.77 0.485 3.835 0.55 ;
      LAYER via2 ;
        RECT 3.7675 0.4825 3.8375 0.5525 ;
    END
  END rd_sel[30]
  PIN rd_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.86 0.45 0.93 0.585 ;
        RECT 0.585 0.9075 0.9275 0.9725 ;
        RECT 0.8625 0.4475 0.9275 0.9725 ;
        RECT 0.215 0.53 0.35 0.595 ;
      LAYER metal2 ;
        RECT 0.86 0.1275 0.93 0.5875 ;
        RECT 0 0.1275 0.93 0.1975 ;
        RECT 0 0.5275 0.35 0.5975 ;
        RECT 0 0.1275 0.07 0.5975 ;
      LAYER metal3 ;
        RECT 0.86 0.055 0.93 1.49 ;
      LAYER via1 ;
        RECT 0.25 0.53 0.315 0.595 ;
        RECT 0.8625 0.485 0.9275 0.55 ;
      LAYER via2 ;
        RECT 0.86 0.4825 0.93 0.5525 ;
    END
  END rd_sel[31]
  PIN rd_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 82.27 0.45 82.34 0.585 ;
        RECT 81.995 0.9075 82.3375 0.9725 ;
        RECT 82.2725 0.4475 82.3375 0.9725 ;
        RECT 81.625 0.53 81.76 0.595 ;
      LAYER metal2 ;
        RECT 82.27 0.12 82.34 0.5875 ;
        RECT 81.41 0.12 82.34 0.19 ;
        RECT 81.41 0.5275 81.76 0.5975 ;
        RECT 81.41 0.12 81.48 0.5975 ;
      LAYER metal3 ;
        RECT 82.27 0.055 82.34 1.4925 ;
      LAYER via1 ;
        RECT 81.66 0.53 81.725 0.595 ;
        RECT 82.2725 0.485 82.3375 0.55 ;
      LAYER via2 ;
        RECT 82.27 0.4825 82.34 0.5525 ;
    END
  END rd_sel[3]
  PIN rd_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 79.3625 0.45 79.4325 0.585 ;
        RECT 79.0875 0.9075 79.43 0.9725 ;
        RECT 79.365 0.4475 79.43 0.9725 ;
        RECT 78.7175 0.53 78.8525 0.595 ;
      LAYER metal2 ;
        RECT 79.3625 0.12 79.4325 0.5875 ;
        RECT 78.5025 0.12 79.4325 0.19 ;
        RECT 78.5025 0.5275 78.8525 0.5975 ;
        RECT 78.5025 0.12 78.5725 0.5975 ;
      LAYER metal3 ;
        RECT 79.3625 0.055 79.4325 1.4925 ;
      LAYER via1 ;
        RECT 78.7525 0.53 78.8175 0.595 ;
        RECT 79.365 0.485 79.43 0.55 ;
      LAYER via2 ;
        RECT 79.3625 0.4825 79.4325 0.5525 ;
    END
  END rd_sel[4]
  PIN rd_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 76.455 0.45 76.525 0.585 ;
        RECT 76.18 0.9075 76.5225 0.9725 ;
        RECT 76.4575 0.4475 76.5225 0.9725 ;
        RECT 75.81 0.53 75.945 0.595 ;
      LAYER metal2 ;
        RECT 76.455 0.12 76.525 0.5875 ;
        RECT 75.595 0.12 76.525 0.19 ;
        RECT 75.595 0.5275 75.945 0.5975 ;
        RECT 75.595 0.12 75.665 0.5975 ;
      LAYER metal3 ;
        RECT 76.455 0.055 76.525 1.4925 ;
      LAYER via1 ;
        RECT 75.845 0.53 75.91 0.595 ;
        RECT 76.4575 0.485 76.5225 0.55 ;
      LAYER via2 ;
        RECT 76.455 0.4825 76.525 0.5525 ;
    END
  END rd_sel[5]
  PIN rd_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 73.5475 0.45 73.6175 0.585 ;
        RECT 73.2725 0.9075 73.615 0.9725 ;
        RECT 73.55 0.4475 73.615 0.9725 ;
        RECT 72.9025 0.53 73.0375 0.595 ;
      LAYER metal2 ;
        RECT 73.5475 0.12 73.6175 0.5875 ;
        RECT 72.6875 0.12 73.6175 0.19 ;
        RECT 72.6875 0.5275 73.0375 0.5975 ;
        RECT 72.6875 0.12 72.7575 0.5975 ;
      LAYER metal3 ;
        RECT 73.5475 0.055 73.6175 1.4925 ;
      LAYER via1 ;
        RECT 72.9375 0.53 73.0025 0.595 ;
        RECT 73.55 0.485 73.615 0.55 ;
      LAYER via2 ;
        RECT 73.5475 0.4825 73.6175 0.5525 ;
    END
  END rd_sel[6]
  PIN rd_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 70.64 0.45 70.71 0.585 ;
        RECT 70.365 0.9075 70.7075 0.9725 ;
        RECT 70.6425 0.4475 70.7075 0.9725 ;
        RECT 69.995 0.53 70.13 0.595 ;
      LAYER metal2 ;
        RECT 70.64 0.12 70.71 0.5875 ;
        RECT 69.78 0.12 70.71 0.19 ;
        RECT 69.78 0.5275 70.13 0.5975 ;
        RECT 69.78 0.12 69.85 0.5975 ;
      LAYER metal3 ;
        RECT 70.64 0.055 70.71 1.4925 ;
      LAYER via1 ;
        RECT 70.03 0.53 70.095 0.595 ;
        RECT 70.6425 0.485 70.7075 0.55 ;
      LAYER via2 ;
        RECT 70.64 0.4825 70.71 0.5525 ;
    END
  END rd_sel[7]
  PIN rd_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 67.7325 0.45 67.8025 0.585 ;
        RECT 67.4575 0.9075 67.8 0.9725 ;
        RECT 67.735 0.4475 67.8 0.9725 ;
        RECT 67.0875 0.53 67.2225 0.595 ;
      LAYER metal2 ;
        RECT 67.7325 0.12 67.8025 0.5875 ;
        RECT 66.8725 0.12 67.8025 0.19 ;
        RECT 66.8725 0.5275 67.2225 0.5975 ;
        RECT 66.8725 0.12 66.9425 0.5975 ;
      LAYER metal3 ;
        RECT 67.7325 0.055 67.8025 1.4925 ;
      LAYER via1 ;
        RECT 67.1225 0.53 67.1875 0.595 ;
        RECT 67.735 0.485 67.8 0.55 ;
      LAYER via2 ;
        RECT 67.7325 0.4825 67.8025 0.5525 ;
    END
  END rd_sel[8]
  PIN rd_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 64.825 0.45 64.895 0.585 ;
        RECT 64.55 0.9075 64.8925 0.9725 ;
        RECT 64.8275 0.4475 64.8925 0.9725 ;
        RECT 64.18 0.53 64.315 0.595 ;
      LAYER metal2 ;
        RECT 64.825 0.12 64.895 0.5875 ;
        RECT 63.965 0.12 64.895 0.19 ;
        RECT 63.965 0.5275 64.315 0.5975 ;
        RECT 63.965 0.12 64.035 0.5975 ;
      LAYER metal3 ;
        RECT 64.825 0.055 64.895 1.4925 ;
      LAYER via1 ;
        RECT 64.215 0.53 64.28 0.595 ;
        RECT 64.8275 0.485 64.8925 0.55 ;
      LAYER via2 ;
        RECT 64.825 0.4825 64.895 0.5525 ;
    END
  END rd_sel[9]
  PIN rd_sel_bar[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 61.6425 0.485 61.7775 0.55 ;
        RECT 61.3975 0.735 61.7425 0.8 ;
        RECT 61.6775 0.485 61.7425 0.8 ;
        RECT 61.3975 0.7 61.4675 0.835 ;
        RECT 61.2725 0.9075 61.465 0.9725 ;
        RECT 61.4 0.675 61.465 0.9725 ;
      LAYER metal2 ;
        RECT 61.3975 0.6975 61.4675 0.8375 ;
      LAYER metal3 ;
        RECT 61.3975 0.055 61.4675 1.4925 ;
      LAYER via1 ;
        RECT 61.4 0.735 61.465 0.8 ;
      LAYER via2 ;
        RECT 61.3975 0.7325 61.4675 0.8025 ;
    END
  END rd_sel_bar[10]
  PIN rd_sel_bar[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 58.735 0.485 58.87 0.55 ;
        RECT 58.49 0.735 58.835 0.8 ;
        RECT 58.77 0.485 58.835 0.8 ;
        RECT 58.49 0.7 58.56 0.835 ;
        RECT 58.365 0.9075 58.5575 0.9725 ;
        RECT 58.4925 0.675 58.5575 0.9725 ;
      LAYER metal2 ;
        RECT 58.49 0.6975 58.56 0.8375 ;
      LAYER metal3 ;
        RECT 58.49 0.055 58.56 1.4925 ;
      LAYER via1 ;
        RECT 58.4925 0.735 58.5575 0.8 ;
      LAYER via2 ;
        RECT 58.49 0.7325 58.56 0.8025 ;
    END
  END rd_sel_bar[11]
  PIN rd_sel_bar[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 55.8275 0.485 55.9625 0.55 ;
        RECT 55.5825 0.735 55.9275 0.8 ;
        RECT 55.8625 0.485 55.9275 0.8 ;
        RECT 55.5825 0.7 55.6525 0.835 ;
        RECT 55.4575 0.9075 55.65 0.9725 ;
        RECT 55.585 0.675 55.65 0.9725 ;
      LAYER metal2 ;
        RECT 55.5825 0.6975 55.6525 0.8375 ;
      LAYER metal3 ;
        RECT 55.5825 0.055 55.6525 1.4925 ;
      LAYER via1 ;
        RECT 55.585 0.735 55.65 0.8 ;
      LAYER via2 ;
        RECT 55.5825 0.7325 55.6525 0.8025 ;
    END
  END rd_sel_bar[12]
  PIN rd_sel_bar[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 52.92 0.485 53.055 0.55 ;
        RECT 52.675 0.735 53.02 0.8 ;
        RECT 52.955 0.485 53.02 0.8 ;
        RECT 52.675 0.7 52.745 0.835 ;
        RECT 52.55 0.9075 52.7425 0.9725 ;
        RECT 52.6775 0.675 52.7425 0.9725 ;
      LAYER metal2 ;
        RECT 52.675 0.6975 52.745 0.8375 ;
      LAYER metal3 ;
        RECT 52.675 0.055 52.745 1.4925 ;
      LAYER via1 ;
        RECT 52.6775 0.735 52.7425 0.8 ;
      LAYER via2 ;
        RECT 52.675 0.7325 52.745 0.8025 ;
    END
  END rd_sel_bar[13]
  PIN rd_sel_bar[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 50.0125 0.485 50.1475 0.55 ;
        RECT 49.7675 0.735 50.1125 0.8 ;
        RECT 50.0475 0.485 50.1125 0.8 ;
        RECT 49.7675 0.7 49.8375 0.835 ;
        RECT 49.6425 0.9075 49.835 0.9725 ;
        RECT 49.77 0.675 49.835 0.9725 ;
      LAYER metal2 ;
        RECT 49.7675 0.6975 49.8375 0.8375 ;
      LAYER metal3 ;
        RECT 49.7675 0.055 49.8375 1.4925 ;
      LAYER via1 ;
        RECT 49.77 0.735 49.835 0.8 ;
      LAYER via2 ;
        RECT 49.7675 0.7325 49.8375 0.8025 ;
    END
  END rd_sel_bar[14]
  PIN rd_sel_bar[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 47.105 0.485 47.24 0.55 ;
        RECT 46.86 0.735 47.205 0.8 ;
        RECT 47.14 0.485 47.205 0.8 ;
        RECT 46.86 0.7 46.93 0.835 ;
        RECT 46.735 0.9075 46.9275 0.9725 ;
        RECT 46.8625 0.675 46.9275 0.9725 ;
      LAYER metal2 ;
        RECT 46.86 0.6975 46.93 0.8375 ;
      LAYER metal3 ;
        RECT 46.86 0.055 46.93 1.4925 ;
      LAYER via1 ;
        RECT 46.8625 0.735 46.9275 0.8 ;
      LAYER via2 ;
        RECT 46.86 0.7325 46.93 0.8025 ;
    END
  END rd_sel_bar[15]
  PIN rd_sel_bar[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 44.1975 0.485 44.3325 0.55 ;
        RECT 43.9525 0.735 44.2975 0.8 ;
        RECT 44.2325 0.485 44.2975 0.8 ;
        RECT 43.9525 0.7 44.0225 0.835 ;
        RECT 43.8275 0.9075 44.02 0.9725 ;
        RECT 43.955 0.675 44.02 0.9725 ;
      LAYER metal2 ;
        RECT 43.9525 0.6975 44.0225 0.8375 ;
      LAYER metal3 ;
        RECT 43.9525 0.055 44.0225 1.4925 ;
      LAYER via1 ;
        RECT 43.955 0.735 44.02 0.8 ;
      LAYER via2 ;
        RECT 43.9525 0.7325 44.0225 0.8025 ;
    END
  END rd_sel_bar[16]
  PIN rd_sel_bar[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 41.29 0.485 41.425 0.55 ;
        RECT 41.045 0.735 41.39 0.8 ;
        RECT 41.325 0.485 41.39 0.8 ;
        RECT 41.045 0.7 41.115 0.835 ;
        RECT 40.92 0.9075 41.1125 0.9725 ;
        RECT 41.0475 0.675 41.1125 0.9725 ;
      LAYER metal2 ;
        RECT 41.045 0.6975 41.115 0.8375 ;
      LAYER metal3 ;
        RECT 41.045 0.055 41.115 1.4925 ;
      LAYER via1 ;
        RECT 41.0475 0.735 41.1125 0.8 ;
      LAYER via2 ;
        RECT 41.045 0.7325 41.115 0.8025 ;
    END
  END rd_sel_bar[17]
  PIN rd_sel_bar[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 38.3825 0.485 38.5175 0.55 ;
        RECT 38.1375 0.735 38.4825 0.8 ;
        RECT 38.4175 0.485 38.4825 0.8 ;
        RECT 38.1375 0.7 38.2075 0.835 ;
        RECT 38.0125 0.9075 38.205 0.9725 ;
        RECT 38.14 0.675 38.205 0.9725 ;
      LAYER metal2 ;
        RECT 38.1375 0.6975 38.2075 0.8375 ;
      LAYER metal3 ;
        RECT 38.1375 0.055 38.2075 1.4925 ;
      LAYER via1 ;
        RECT 38.14 0.735 38.205 0.8 ;
      LAYER via2 ;
        RECT 38.1375 0.7325 38.2075 0.8025 ;
    END
  END rd_sel_bar[18]
  PIN rd_sel_bar[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 35.475 0.485 35.61 0.55 ;
        RECT 35.23 0.735 35.575 0.8 ;
        RECT 35.51 0.485 35.575 0.8 ;
        RECT 35.23 0.7 35.3 0.835 ;
        RECT 35.105 0.9075 35.2975 0.9725 ;
        RECT 35.2325 0.675 35.2975 0.9725 ;
      LAYER metal2 ;
        RECT 35.23 0.6975 35.3 0.8375 ;
      LAYER metal3 ;
        RECT 35.23 0.055 35.3 1.4925 ;
      LAYER via1 ;
        RECT 35.2325 0.735 35.2975 0.8 ;
      LAYER via2 ;
        RECT 35.23 0.7325 35.3 0.8025 ;
    END
  END rd_sel_bar[19]
  PIN rd_sel_bar[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 87.81 0.485 87.945 0.55 ;
        RECT 87.565 0.735 87.91 0.8 ;
        RECT 87.845 0.485 87.91 0.8 ;
        RECT 87.565 0.7 87.635 0.835 ;
        RECT 87.44 0.9075 87.6325 0.9725 ;
        RECT 87.5675 0.675 87.6325 0.9725 ;
      LAYER metal2 ;
        RECT 87.565 0.6975 87.635 0.8375 ;
      LAYER metal3 ;
        RECT 87.565 0.055 87.635 1.4925 ;
      LAYER via1 ;
        RECT 87.5675 0.735 87.6325 0.8 ;
      LAYER via2 ;
        RECT 87.565 0.7325 87.635 0.8025 ;
    END
  END rd_sel_bar[1]
  PIN rd_sel_bar[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 32.5675 0.485 32.7025 0.55 ;
        RECT 32.3225 0.735 32.6675 0.8 ;
        RECT 32.6025 0.485 32.6675 0.8 ;
        RECT 32.3225 0.7 32.3925 0.835 ;
        RECT 32.1975 0.9075 32.39 0.9725 ;
        RECT 32.325 0.675 32.39 0.9725 ;
      LAYER metal2 ;
        RECT 32.3225 0.6975 32.3925 0.8375 ;
      LAYER metal3 ;
        RECT 32.3225 0.055 32.3925 1.4925 ;
      LAYER via1 ;
        RECT 32.325 0.735 32.39 0.8 ;
      LAYER via2 ;
        RECT 32.3225 0.7325 32.3925 0.8025 ;
    END
  END rd_sel_bar[20]
  PIN rd_sel_bar[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 29.66 0.485 29.795 0.55 ;
        RECT 29.415 0.735 29.76 0.8 ;
        RECT 29.695 0.485 29.76 0.8 ;
        RECT 29.415 0.7 29.485 0.835 ;
        RECT 29.29 0.9075 29.4825 0.9725 ;
        RECT 29.4175 0.675 29.4825 0.9725 ;
      LAYER metal2 ;
        RECT 29.415 0.6975 29.485 0.8375 ;
      LAYER metal3 ;
        RECT 29.415 0.055 29.485 1.4925 ;
      LAYER via1 ;
        RECT 29.4175 0.735 29.4825 0.8 ;
      LAYER via2 ;
        RECT 29.415 0.7325 29.485 0.8025 ;
    END
  END rd_sel_bar[21]
  PIN rd_sel_bar[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 26.7525 0.485 26.8875 0.55 ;
        RECT 26.5075 0.735 26.8525 0.8 ;
        RECT 26.7875 0.485 26.8525 0.8 ;
        RECT 26.5075 0.7 26.5775 0.835 ;
        RECT 26.3825 0.9075 26.575 0.9725 ;
        RECT 26.51 0.675 26.575 0.9725 ;
      LAYER metal2 ;
        RECT 26.5075 0.6975 26.5775 0.8375 ;
      LAYER metal3 ;
        RECT 26.5075 0.055 26.5775 1.4925 ;
      LAYER via1 ;
        RECT 26.51 0.735 26.575 0.8 ;
      LAYER via2 ;
        RECT 26.5075 0.7325 26.5775 0.8025 ;
    END
  END rd_sel_bar[22]
  PIN rd_sel_bar[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 23.845 0.485 23.98 0.55 ;
        RECT 23.6 0.735 23.945 0.8 ;
        RECT 23.88 0.485 23.945 0.8 ;
        RECT 23.6 0.7 23.67 0.835 ;
        RECT 23.475 0.9075 23.6675 0.9725 ;
        RECT 23.6025 0.675 23.6675 0.9725 ;
      LAYER metal2 ;
        RECT 23.6 0.6975 23.67 0.8375 ;
      LAYER metal3 ;
        RECT 23.6 0.055 23.67 1.4925 ;
      LAYER via1 ;
        RECT 23.6025 0.735 23.6675 0.8 ;
      LAYER via2 ;
        RECT 23.6 0.7325 23.67 0.8025 ;
    END
  END rd_sel_bar[23]
  PIN rd_sel_bar[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 20.9375 0.485 21.0725 0.55 ;
        RECT 20.6925 0.735 21.0375 0.8 ;
        RECT 20.9725 0.485 21.0375 0.8 ;
        RECT 20.6925 0.7 20.7625 0.835 ;
        RECT 20.5675 0.9075 20.76 0.9725 ;
        RECT 20.695 0.675 20.76 0.9725 ;
      LAYER metal2 ;
        RECT 20.6925 0.6975 20.7625 0.8375 ;
      LAYER metal3 ;
        RECT 20.6925 0.055 20.7625 1.4925 ;
      LAYER via1 ;
        RECT 20.695 0.735 20.76 0.8 ;
      LAYER via2 ;
        RECT 20.6925 0.7325 20.7625 0.8025 ;
    END
  END rd_sel_bar[24]
  PIN rd_sel_bar[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 18.03 0.485 18.165 0.55 ;
        RECT 17.785 0.735 18.13 0.8 ;
        RECT 18.065 0.485 18.13 0.8 ;
        RECT 17.785 0.7 17.855 0.835 ;
        RECT 17.66 0.9075 17.8525 0.9725 ;
        RECT 17.7875 0.675 17.8525 0.9725 ;
      LAYER metal2 ;
        RECT 17.785 0.6975 17.855 0.8375 ;
      LAYER metal3 ;
        RECT 17.785 0.055 17.855 1.4925 ;
      LAYER via1 ;
        RECT 17.7875 0.735 17.8525 0.8 ;
      LAYER via2 ;
        RECT 17.785 0.7325 17.855 0.8025 ;
    END
  END rd_sel_bar[25]
  PIN rd_sel_bar[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.1225 0.485 15.2575 0.55 ;
        RECT 14.8775 0.735 15.2225 0.8 ;
        RECT 15.1575 0.485 15.2225 0.8 ;
        RECT 14.8775 0.7 14.9475 0.835 ;
        RECT 14.7525 0.9075 14.945 0.9725 ;
        RECT 14.88 0.675 14.945 0.9725 ;
      LAYER metal2 ;
        RECT 14.8775 0.6975 14.9475 0.8375 ;
      LAYER metal3 ;
        RECT 14.8775 0.055 14.9475 1.4925 ;
      LAYER via1 ;
        RECT 14.88 0.735 14.945 0.8 ;
      LAYER via2 ;
        RECT 14.8775 0.7325 14.9475 0.8025 ;
    END
  END rd_sel_bar[26]
  PIN rd_sel_bar[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.215 0.485 12.35 0.55 ;
        RECT 11.97 0.735 12.315 0.8 ;
        RECT 12.25 0.485 12.315 0.8 ;
        RECT 11.97 0.7 12.04 0.835 ;
        RECT 11.845 0.9075 12.0375 0.9725 ;
        RECT 11.9725 0.675 12.0375 0.9725 ;
      LAYER metal2 ;
        RECT 11.97 0.6975 12.04 0.8375 ;
      LAYER metal3 ;
        RECT 11.97 0.055 12.04 1.4925 ;
      LAYER via1 ;
        RECT 11.9725 0.735 12.0375 0.8 ;
      LAYER via2 ;
        RECT 11.97 0.7325 12.04 0.8025 ;
    END
  END rd_sel_bar[27]
  PIN rd_sel_bar[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.3075 0.485 9.4425 0.55 ;
        RECT 9.0625 0.735 9.4075 0.8 ;
        RECT 9.3425 0.485 9.4075 0.8 ;
        RECT 9.0625 0.7 9.1325 0.835 ;
        RECT 8.9375 0.9075 9.13 0.9725 ;
        RECT 9.065 0.675 9.13 0.9725 ;
      LAYER metal2 ;
        RECT 9.0625 0.6975 9.1325 0.8375 ;
      LAYER metal3 ;
        RECT 9.0625 0.055 9.1325 1.4925 ;
      LAYER via1 ;
        RECT 9.065 0.735 9.13 0.8 ;
      LAYER via2 ;
        RECT 9.0625 0.7325 9.1325 0.8025 ;
    END
  END rd_sel_bar[28]
  PIN rd_sel_bar[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.4 0.485 6.535 0.55 ;
        RECT 6.155 0.735 6.5 0.8 ;
        RECT 6.435 0.485 6.5 0.8 ;
        RECT 6.155 0.7 6.225 0.835 ;
        RECT 6.03 0.9075 6.2225 0.9725 ;
        RECT 6.1575 0.675 6.2225 0.9725 ;
      LAYER metal2 ;
        RECT 6.155 0.6975 6.225 0.8375 ;
      LAYER metal3 ;
        RECT 6.155 0.055 6.225 1.4925 ;
      LAYER via1 ;
        RECT 6.1575 0.735 6.2225 0.8 ;
      LAYER via2 ;
        RECT 6.155 0.7325 6.225 0.8025 ;
    END
  END rd_sel_bar[29]
  PIN rd_sel_bar[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 84.9025 0.485 85.0375 0.55 ;
        RECT 84.6575 0.735 85.0025 0.8 ;
        RECT 84.9375 0.485 85.0025 0.8 ;
        RECT 84.6575 0.7 84.7275 0.835 ;
        RECT 84.5325 0.9075 84.725 0.9725 ;
        RECT 84.66 0.675 84.725 0.9725 ;
      LAYER metal2 ;
        RECT 84.6575 0.6975 84.7275 0.8375 ;
      LAYER metal3 ;
        RECT 84.6575 0.055 84.7275 1.4925 ;
      LAYER via1 ;
        RECT 84.66 0.735 84.725 0.8 ;
      LAYER via2 ;
        RECT 84.6575 0.7325 84.7275 0.8025 ;
    END
  END rd_sel_bar[2]
  PIN rd_sel_bar[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.4925 0.485 3.6275 0.55 ;
        RECT 3.2475 0.735 3.5925 0.8 ;
        RECT 3.5275 0.485 3.5925 0.8 ;
        RECT 3.2475 0.7 3.3175 0.835 ;
        RECT 3.1225 0.9075 3.315 0.9725 ;
        RECT 3.25 0.675 3.315 0.9725 ;
      LAYER metal2 ;
        RECT 3.2475 0.6975 3.3175 0.8375 ;
      LAYER metal3 ;
        RECT 3.2475 0.055 3.3175 1.4925 ;
      LAYER via1 ;
        RECT 3.25 0.735 3.315 0.8 ;
      LAYER via2 ;
        RECT 3.2475 0.7325 3.3175 0.8025 ;
    END
  END rd_sel_bar[30]
  PIN rd_sel_bar[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.585 0.485 0.72 0.55 ;
        RECT 0.34 0.735 0.685 0.8 ;
        RECT 0.62 0.485 0.685 0.8 ;
        RECT 0.34 0.7 0.41 0.835 ;
        RECT 0.215 0.9075 0.4075 0.9725 ;
        RECT 0.3425 0.675 0.4075 0.9725 ;
      LAYER metal2 ;
        RECT 0.34 0.6975 0.41 0.8375 ;
      LAYER metal3 ;
        RECT 0.34 0.055 0.41 1.49 ;
      LAYER via1 ;
        RECT 0.3425 0.735 0.4075 0.8 ;
      LAYER via2 ;
        RECT 0.34 0.7325 0.41 0.8025 ;
    END
  END rd_sel_bar[31]
  PIN rd_sel_bar[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 81.995 0.485 82.13 0.55 ;
        RECT 81.75 0.735 82.095 0.8 ;
        RECT 82.03 0.485 82.095 0.8 ;
        RECT 81.75 0.7 81.82 0.835 ;
        RECT 81.625 0.9075 81.8175 0.9725 ;
        RECT 81.7525 0.675 81.8175 0.9725 ;
      LAYER metal2 ;
        RECT 81.75 0.6975 81.82 0.8375 ;
      LAYER metal3 ;
        RECT 81.75 0.055 81.82 1.4925 ;
      LAYER via1 ;
        RECT 81.7525 0.735 81.8175 0.8 ;
      LAYER via2 ;
        RECT 81.75 0.7325 81.82 0.8025 ;
    END
  END rd_sel_bar[3]
  PIN rd_sel_bar[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 79.0875 0.485 79.2225 0.55 ;
        RECT 78.8425 0.735 79.1875 0.8 ;
        RECT 79.1225 0.485 79.1875 0.8 ;
        RECT 78.8425 0.7 78.9125 0.835 ;
        RECT 78.7175 0.9075 78.91 0.9725 ;
        RECT 78.845 0.675 78.91 0.9725 ;
      LAYER metal2 ;
        RECT 78.8425 0.6975 78.9125 0.8375 ;
      LAYER metal3 ;
        RECT 78.8425 0.055 78.9125 1.4925 ;
      LAYER via1 ;
        RECT 78.845 0.735 78.91 0.8 ;
      LAYER via2 ;
        RECT 78.8425 0.7325 78.9125 0.8025 ;
    END
  END rd_sel_bar[4]
  PIN rd_sel_bar[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 76.18 0.485 76.315 0.55 ;
        RECT 75.935 0.735 76.28 0.8 ;
        RECT 76.215 0.485 76.28 0.8 ;
        RECT 75.935 0.7 76.005 0.835 ;
        RECT 75.81 0.9075 76.0025 0.9725 ;
        RECT 75.9375 0.675 76.0025 0.9725 ;
      LAYER metal2 ;
        RECT 75.935 0.6975 76.005 0.8375 ;
      LAYER metal3 ;
        RECT 75.935 0.055 76.005 1.4925 ;
      LAYER via1 ;
        RECT 75.9375 0.735 76.0025 0.8 ;
      LAYER via2 ;
        RECT 75.935 0.7325 76.005 0.8025 ;
    END
  END rd_sel_bar[5]
  PIN rd_sel_bar[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 73.2725 0.485 73.4075 0.55 ;
        RECT 73.0275 0.735 73.3725 0.8 ;
        RECT 73.3075 0.485 73.3725 0.8 ;
        RECT 73.0275 0.7 73.0975 0.835 ;
        RECT 72.9025 0.9075 73.095 0.9725 ;
        RECT 73.03 0.675 73.095 0.9725 ;
      LAYER metal2 ;
        RECT 73.0275 0.6975 73.0975 0.8375 ;
      LAYER metal3 ;
        RECT 73.0275 0.055 73.0975 1.4925 ;
      LAYER via1 ;
        RECT 73.03 0.735 73.095 0.8 ;
      LAYER via2 ;
        RECT 73.0275 0.7325 73.0975 0.8025 ;
    END
  END rd_sel_bar[6]
  PIN rd_sel_bar[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 70.365 0.485 70.5 0.55 ;
        RECT 70.12 0.735 70.465 0.8 ;
        RECT 70.4 0.485 70.465 0.8 ;
        RECT 70.12 0.7 70.19 0.835 ;
        RECT 69.995 0.9075 70.1875 0.9725 ;
        RECT 70.1225 0.675 70.1875 0.9725 ;
      LAYER metal2 ;
        RECT 70.12 0.6975 70.19 0.8375 ;
      LAYER metal3 ;
        RECT 70.12 0.055 70.19 1.4925 ;
      LAYER via1 ;
        RECT 70.1225 0.735 70.1875 0.8 ;
      LAYER via2 ;
        RECT 70.12 0.7325 70.19 0.8025 ;
    END
  END rd_sel_bar[7]
  PIN rd_sel_bar[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 67.4575 0.485 67.5925 0.55 ;
        RECT 67.2125 0.735 67.5575 0.8 ;
        RECT 67.4925 0.485 67.5575 0.8 ;
        RECT 67.2125 0.7 67.2825 0.835 ;
        RECT 67.0875 0.9075 67.28 0.9725 ;
        RECT 67.215 0.675 67.28 0.9725 ;
      LAYER metal2 ;
        RECT 67.2125 0.6975 67.2825 0.8375 ;
      LAYER metal3 ;
        RECT 67.2125 0.055 67.2825 1.4925 ;
      LAYER via1 ;
        RECT 67.215 0.735 67.28 0.8 ;
      LAYER via2 ;
        RECT 67.2125 0.7325 67.2825 0.8025 ;
    END
  END rd_sel_bar[8]
  PIN rd_sel_bar[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 64.55 0.485 64.685 0.55 ;
        RECT 64.305 0.735 64.65 0.8 ;
        RECT 64.585 0.485 64.65 0.8 ;
        RECT 64.305 0.7 64.375 0.835 ;
        RECT 64.18 0.9075 64.3725 0.9725 ;
        RECT 64.3075 0.675 64.3725 0.9725 ;
      LAYER metal2 ;
        RECT 64.305 0.6975 64.375 0.8375 ;
      LAYER metal3 ;
        RECT 64.305 0.055 64.375 1.4925 ;
      LAYER via1 ;
        RECT 64.3075 0.735 64.3725 0.8 ;
      LAYER via2 ;
        RECT 64.305 0.7325 64.375 0.8025 ;
    END
  END rd_sel_bar[9]
  PIN rs1_rdata
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 93.645 0.5825 93.715 0.7175 ;
        RECT 93.645 0.265 93.71 1.285 ;
        RECT 93.39 0.5325 93.71 0.5975 ;
        RECT 93.39 0.4975 93.455 0.6325 ;
      LAYER metal2 ;
        RECT 93.645 0.58 93.715 0.72 ;
      LAYER metal3 ;
        RECT 93.645 0.055 93.715 1.4925 ;
      LAYER via1 ;
        RECT 93.6475 0.6175 93.7125 0.6825 ;
      LAYER via2 ;
        RECT 93.645 0.615 93.715 0.685 ;
    END
  END rs1_rdata
  PIN rs1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 91.6475 0.785 91.7175 0.92 ;
        RECT 91.3675 0.485 91.7175 0.55 ;
        RECT 91.65 0.4825 91.715 0.9225 ;
      LAYER metal2 ;
        RECT 91.6475 0.7825 91.7175 0.9225 ;
      LAYER metal3 ;
        RECT 91.6475 0.055 91.7175 1.4925 ;
      LAYER via1 ;
        RECT 91.65 0.82 91.715 0.885 ;
      LAYER via2 ;
        RECT 91.6475 0.8175 91.7175 0.8875 ;
    END
  END rs1_sel[0]
  PIN rs1_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.8725 0.785 63.9425 0.92 ;
        RECT 63.5925 0.485 63.9425 0.55 ;
        RECT 63.875 0.4825 63.94 0.9225 ;
      LAYER metal2 ;
        RECT 63.8725 0.7825 63.9425 0.9225 ;
      LAYER metal3 ;
        RECT 63.8725 0.055 63.9425 1.4925 ;
      LAYER via1 ;
        RECT 63.875 0.82 63.94 0.885 ;
      LAYER via2 ;
        RECT 63.8725 0.8175 63.9425 0.8875 ;
    END
  END rs1_sel[10]
  PIN rs1_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 60.965 0.785 61.035 0.92 ;
        RECT 60.685 0.485 61.035 0.55 ;
        RECT 60.9675 0.4825 61.0325 0.9225 ;
      LAYER metal2 ;
        RECT 60.965 0.7825 61.035 0.9225 ;
      LAYER metal3 ;
        RECT 60.965 0.055 61.035 1.4925 ;
      LAYER via1 ;
        RECT 60.9675 0.82 61.0325 0.885 ;
      LAYER via2 ;
        RECT 60.965 0.8175 61.035 0.8875 ;
    END
  END rs1_sel[11]
  PIN rs1_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 58.0575 0.785 58.1275 0.92 ;
        RECT 57.7775 0.485 58.1275 0.55 ;
        RECT 58.06 0.4825 58.125 0.9225 ;
      LAYER metal2 ;
        RECT 58.0575 0.7825 58.1275 0.9225 ;
      LAYER metal3 ;
        RECT 58.0575 0.055 58.1275 1.4925 ;
      LAYER via1 ;
        RECT 58.06 0.82 58.125 0.885 ;
      LAYER via2 ;
        RECT 58.0575 0.8175 58.1275 0.8875 ;
    END
  END rs1_sel[12]
  PIN rs1_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 55.15 0.785 55.22 0.92 ;
        RECT 54.87 0.485 55.22 0.55 ;
        RECT 55.1525 0.4825 55.2175 0.9225 ;
      LAYER metal2 ;
        RECT 55.15 0.7825 55.22 0.9225 ;
      LAYER metal3 ;
        RECT 55.15 0.055 55.22 1.4925 ;
      LAYER via1 ;
        RECT 55.1525 0.82 55.2175 0.885 ;
      LAYER via2 ;
        RECT 55.15 0.8175 55.22 0.8875 ;
    END
  END rs1_sel[13]
  PIN rs1_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 52.2425 0.785 52.3125 0.92 ;
        RECT 51.9625 0.485 52.3125 0.55 ;
        RECT 52.245 0.4825 52.31 0.9225 ;
      LAYER metal2 ;
        RECT 52.2425 0.7825 52.3125 0.9225 ;
      LAYER metal3 ;
        RECT 52.2425 0.055 52.3125 1.4925 ;
      LAYER via1 ;
        RECT 52.245 0.82 52.31 0.885 ;
      LAYER via2 ;
        RECT 52.2425 0.8175 52.3125 0.8875 ;
    END
  END rs1_sel[14]
  PIN rs1_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 49.335 0.785 49.405 0.92 ;
        RECT 49.055 0.485 49.405 0.55 ;
        RECT 49.3375 0.4825 49.4025 0.9225 ;
      LAYER metal2 ;
        RECT 49.335 0.7825 49.405 0.9225 ;
      LAYER metal3 ;
        RECT 49.335 0.055 49.405 1.4925 ;
      LAYER via1 ;
        RECT 49.3375 0.82 49.4025 0.885 ;
      LAYER via2 ;
        RECT 49.335 0.8175 49.405 0.8875 ;
    END
  END rs1_sel[15]
  PIN rs1_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 46.4275 0.785 46.4975 0.92 ;
        RECT 46.1475 0.485 46.4975 0.55 ;
        RECT 46.43 0.4825 46.495 0.9225 ;
      LAYER metal2 ;
        RECT 46.4275 0.7825 46.4975 0.9225 ;
      LAYER metal3 ;
        RECT 46.4275 0.055 46.4975 1.4925 ;
      LAYER via1 ;
        RECT 46.43 0.82 46.495 0.885 ;
      LAYER via2 ;
        RECT 46.4275 0.8175 46.4975 0.8875 ;
    END
  END rs1_sel[16]
  PIN rs1_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 43.52 0.785 43.59 0.92 ;
        RECT 43.24 0.485 43.59 0.55 ;
        RECT 43.5225 0.4825 43.5875 0.9225 ;
      LAYER metal2 ;
        RECT 43.52 0.7825 43.59 0.9225 ;
      LAYER metal3 ;
        RECT 43.52 0.055 43.59 1.4925 ;
      LAYER via1 ;
        RECT 43.5225 0.82 43.5875 0.885 ;
      LAYER via2 ;
        RECT 43.52 0.8175 43.59 0.8875 ;
    END
  END rs1_sel[17]
  PIN rs1_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 40.6125 0.785 40.6825 0.92 ;
        RECT 40.3325 0.485 40.6825 0.55 ;
        RECT 40.615 0.4825 40.68 0.9225 ;
      LAYER metal2 ;
        RECT 40.6125 0.7825 40.6825 0.9225 ;
      LAYER metal3 ;
        RECT 40.6125 0.055 40.6825 1.4925 ;
      LAYER via1 ;
        RECT 40.615 0.82 40.68 0.885 ;
      LAYER via2 ;
        RECT 40.6125 0.8175 40.6825 0.8875 ;
    END
  END rs1_sel[18]
  PIN rs1_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 37.705 0.785 37.775 0.92 ;
        RECT 37.425 0.485 37.775 0.55 ;
        RECT 37.7075 0.4825 37.7725 0.9225 ;
      LAYER metal2 ;
        RECT 37.705 0.7825 37.775 0.9225 ;
      LAYER metal3 ;
        RECT 37.705 0.055 37.775 1.4925 ;
      LAYER via1 ;
        RECT 37.7075 0.82 37.7725 0.885 ;
      LAYER via2 ;
        RECT 37.705 0.8175 37.775 0.8875 ;
    END
  END rs1_sel[19]
  PIN rs1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 90.04 0.785 90.11 0.92 ;
        RECT 89.76 0.485 90.11 0.55 ;
        RECT 90.0425 0.4825 90.1075 0.9225 ;
      LAYER metal2 ;
        RECT 90.04 0.7825 90.11 0.9225 ;
      LAYER metal3 ;
        RECT 90.04 0.055 90.11 1.4925 ;
      LAYER via1 ;
        RECT 90.0425 0.82 90.1075 0.885 ;
      LAYER via2 ;
        RECT 90.04 0.8175 90.11 0.8875 ;
    END
  END rs1_sel[1]
  PIN rs1_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 34.7975 0.785 34.8675 0.92 ;
        RECT 34.5175 0.485 34.8675 0.55 ;
        RECT 34.8 0.4825 34.865 0.9225 ;
      LAYER metal2 ;
        RECT 34.7975 0.7825 34.8675 0.9225 ;
      LAYER metal3 ;
        RECT 34.7975 0.055 34.8675 1.4925 ;
      LAYER via1 ;
        RECT 34.8 0.82 34.865 0.885 ;
      LAYER via2 ;
        RECT 34.7975 0.8175 34.8675 0.8875 ;
    END
  END rs1_sel[20]
  PIN rs1_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 31.89 0.785 31.96 0.92 ;
        RECT 31.61 0.485 31.96 0.55 ;
        RECT 31.8925 0.4825 31.9575 0.9225 ;
      LAYER metal2 ;
        RECT 31.89 0.7825 31.96 0.9225 ;
      LAYER metal3 ;
        RECT 31.89 0.055 31.96 1.4925 ;
      LAYER via1 ;
        RECT 31.8925 0.82 31.9575 0.885 ;
      LAYER via2 ;
        RECT 31.89 0.8175 31.96 0.8875 ;
    END
  END rs1_sel[21]
  PIN rs1_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 28.9825 0.785 29.0525 0.92 ;
        RECT 28.7025 0.485 29.0525 0.55 ;
        RECT 28.985 0.4825 29.05 0.9225 ;
      LAYER metal2 ;
        RECT 28.9825 0.7825 29.0525 0.9225 ;
      LAYER metal3 ;
        RECT 28.9825 0.055 29.0525 1.4925 ;
      LAYER via1 ;
        RECT 28.985 0.82 29.05 0.885 ;
      LAYER via2 ;
        RECT 28.9825 0.8175 29.0525 0.8875 ;
    END
  END rs1_sel[22]
  PIN rs1_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 26.075 0.785 26.145 0.92 ;
        RECT 25.795 0.485 26.145 0.55 ;
        RECT 26.0775 0.4825 26.1425 0.9225 ;
      LAYER metal2 ;
        RECT 26.075 0.7825 26.145 0.9225 ;
      LAYER metal3 ;
        RECT 26.075 0.055 26.145 1.4925 ;
      LAYER via1 ;
        RECT 26.0775 0.82 26.1425 0.885 ;
      LAYER via2 ;
        RECT 26.075 0.8175 26.145 0.8875 ;
    END
  END rs1_sel[23]
  PIN rs1_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 23.1675 0.785 23.2375 0.92 ;
        RECT 22.8875 0.485 23.2375 0.55 ;
        RECT 23.17 0.4825 23.235 0.9225 ;
      LAYER metal2 ;
        RECT 23.1675 0.7825 23.2375 0.9225 ;
      LAYER metal3 ;
        RECT 23.1675 0.055 23.2375 1.4925 ;
      LAYER via1 ;
        RECT 23.17 0.82 23.235 0.885 ;
      LAYER via2 ;
        RECT 23.1675 0.8175 23.2375 0.8875 ;
    END
  END rs1_sel[24]
  PIN rs1_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 20.26 0.785 20.33 0.92 ;
        RECT 19.98 0.485 20.33 0.55 ;
        RECT 20.2625 0.4825 20.3275 0.9225 ;
      LAYER metal2 ;
        RECT 20.26 0.7825 20.33 0.9225 ;
      LAYER metal3 ;
        RECT 20.26 0.055 20.33 1.4925 ;
      LAYER via1 ;
        RECT 20.2625 0.82 20.3275 0.885 ;
      LAYER via2 ;
        RECT 20.26 0.8175 20.33 0.8875 ;
    END
  END rs1_sel[25]
  PIN rs1_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 17.3525 0.785 17.4225 0.92 ;
        RECT 17.0725 0.485 17.4225 0.55 ;
        RECT 17.355 0.4825 17.42 0.9225 ;
      LAYER metal2 ;
        RECT 17.3525 0.7825 17.4225 0.9225 ;
      LAYER metal3 ;
        RECT 17.3525 0.055 17.4225 1.4925 ;
      LAYER via1 ;
        RECT 17.355 0.82 17.42 0.885 ;
      LAYER via2 ;
        RECT 17.3525 0.8175 17.4225 0.8875 ;
    END
  END rs1_sel[26]
  PIN rs1_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 14.445 0.785 14.515 0.92 ;
        RECT 14.165 0.485 14.515 0.55 ;
        RECT 14.4475 0.4825 14.5125 0.9225 ;
      LAYER metal2 ;
        RECT 14.445 0.7825 14.515 0.9225 ;
      LAYER metal3 ;
        RECT 14.445 0.055 14.515 1.4925 ;
      LAYER via1 ;
        RECT 14.4475 0.82 14.5125 0.885 ;
      LAYER via2 ;
        RECT 14.445 0.8175 14.515 0.8875 ;
    END
  END rs1_sel[27]
  PIN rs1_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 11.5375 0.785 11.6075 0.92 ;
        RECT 11.2575 0.485 11.6075 0.55 ;
        RECT 11.54 0.4825 11.605 0.9225 ;
      LAYER metal2 ;
        RECT 11.5375 0.7825 11.6075 0.9225 ;
      LAYER metal3 ;
        RECT 11.5375 0.055 11.6075 1.4925 ;
      LAYER via1 ;
        RECT 11.54 0.82 11.605 0.885 ;
      LAYER via2 ;
        RECT 11.5375 0.8175 11.6075 0.8875 ;
    END
  END rs1_sel[28]
  PIN rs1_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 8.63 0.785 8.7 0.92 ;
        RECT 8.35 0.485 8.7 0.55 ;
        RECT 8.6325 0.4825 8.6975 0.9225 ;
      LAYER metal2 ;
        RECT 8.63 0.7825 8.7 0.9225 ;
      LAYER metal3 ;
        RECT 8.63 0.055 8.7 1.4925 ;
      LAYER via1 ;
        RECT 8.6325 0.82 8.6975 0.885 ;
      LAYER via2 ;
        RECT 8.63 0.8175 8.7 0.8875 ;
    END
  END rs1_sel[29]
  PIN rs1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 87.1325 0.785 87.2025 0.92 ;
        RECT 86.8525 0.485 87.2025 0.55 ;
        RECT 87.135 0.4825 87.2 0.9225 ;
      LAYER metal2 ;
        RECT 87.1325 0.7825 87.2025 0.9225 ;
      LAYER metal3 ;
        RECT 87.1325 0.055 87.2025 1.4925 ;
      LAYER via1 ;
        RECT 87.135 0.82 87.2 0.885 ;
      LAYER via2 ;
        RECT 87.1325 0.8175 87.2025 0.8875 ;
    END
  END rs1_sel[2]
  PIN rs1_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.7225 0.785 5.7925 0.92 ;
        RECT 5.4425 0.485 5.7925 0.55 ;
        RECT 5.725 0.4825 5.79 0.9225 ;
      LAYER metal2 ;
        RECT 5.7225 0.7825 5.7925 0.9225 ;
      LAYER metal3 ;
        RECT 5.7225 0.055 5.7925 1.4925 ;
      LAYER via1 ;
        RECT 5.725 0.82 5.79 0.885 ;
      LAYER via2 ;
        RECT 5.7225 0.8175 5.7925 0.8875 ;
    END
  END rs1_sel[30]
  PIN rs1_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.815 0.785 2.885 0.92 ;
        RECT 2.535 0.485 2.885 0.55 ;
        RECT 2.8175 0.4825 2.8825 0.9225 ;
      LAYER metal2 ;
        RECT 2.815 0.7825 2.885 0.9225 ;
      LAYER metal3 ;
        RECT 2.815 0.055 2.885 1.49 ;
      LAYER via1 ;
        RECT 2.8175 0.82 2.8825 0.885 ;
      LAYER via2 ;
        RECT 2.815 0.8175 2.885 0.8875 ;
    END
  END rs1_sel[31]
  PIN rs1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 84.225 0.785 84.295 0.92 ;
        RECT 83.945 0.485 84.295 0.55 ;
        RECT 84.2275 0.4825 84.2925 0.9225 ;
      LAYER metal2 ;
        RECT 84.225 0.7825 84.295 0.9225 ;
      LAYER metal3 ;
        RECT 84.225 0.055 84.295 1.4925 ;
      LAYER via1 ;
        RECT 84.2275 0.82 84.2925 0.885 ;
      LAYER via2 ;
        RECT 84.225 0.8175 84.295 0.8875 ;
    END
  END rs1_sel[3]
  PIN rs1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 81.3175 0.785 81.3875 0.92 ;
        RECT 81.0375 0.485 81.3875 0.55 ;
        RECT 81.32 0.4825 81.385 0.9225 ;
      LAYER metal2 ;
        RECT 81.3175 0.7825 81.3875 0.9225 ;
      LAYER metal3 ;
        RECT 81.3175 0.055 81.3875 1.4925 ;
      LAYER via1 ;
        RECT 81.32 0.82 81.385 0.885 ;
      LAYER via2 ;
        RECT 81.3175 0.8175 81.3875 0.8875 ;
    END
  END rs1_sel[4]
  PIN rs1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 78.41 0.785 78.48 0.92 ;
        RECT 78.13 0.485 78.48 0.55 ;
        RECT 78.4125 0.4825 78.4775 0.9225 ;
      LAYER metal2 ;
        RECT 78.41 0.7825 78.48 0.9225 ;
      LAYER metal3 ;
        RECT 78.41 0.055 78.48 1.4925 ;
      LAYER via1 ;
        RECT 78.4125 0.82 78.4775 0.885 ;
      LAYER via2 ;
        RECT 78.41 0.8175 78.48 0.8875 ;
    END
  END rs1_sel[5]
  PIN rs1_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 75.5025 0.785 75.5725 0.92 ;
        RECT 75.2225 0.485 75.5725 0.55 ;
        RECT 75.505 0.4825 75.57 0.9225 ;
      LAYER metal2 ;
        RECT 75.5025 0.7825 75.5725 0.9225 ;
      LAYER metal3 ;
        RECT 75.5025 0.055 75.5725 1.4925 ;
      LAYER via1 ;
        RECT 75.505 0.82 75.57 0.885 ;
      LAYER via2 ;
        RECT 75.5025 0.8175 75.5725 0.8875 ;
    END
  END rs1_sel[6]
  PIN rs1_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 72.595 0.785 72.665 0.92 ;
        RECT 72.315 0.485 72.665 0.55 ;
        RECT 72.5975 0.4825 72.6625 0.9225 ;
      LAYER metal2 ;
        RECT 72.595 0.7825 72.665 0.9225 ;
      LAYER metal3 ;
        RECT 72.595 0.055 72.665 1.4925 ;
      LAYER via1 ;
        RECT 72.5975 0.82 72.6625 0.885 ;
      LAYER via2 ;
        RECT 72.595 0.8175 72.665 0.8875 ;
    END
  END rs1_sel[7]
  PIN rs1_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 69.6875 0.785 69.7575 0.92 ;
        RECT 69.4075 0.485 69.7575 0.55 ;
        RECT 69.69 0.4825 69.755 0.9225 ;
      LAYER metal2 ;
        RECT 69.6875 0.7825 69.7575 0.9225 ;
      LAYER metal3 ;
        RECT 69.6875 0.055 69.7575 1.4925 ;
      LAYER via1 ;
        RECT 69.69 0.82 69.755 0.885 ;
      LAYER via2 ;
        RECT 69.6875 0.8175 69.7575 0.8875 ;
    END
  END rs1_sel[8]
  PIN rs1_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 66.78 0.785 66.85 0.92 ;
        RECT 66.5 0.485 66.85 0.55 ;
        RECT 66.7825 0.4825 66.8475 0.9225 ;
      LAYER metal2 ;
        RECT 66.78 0.7825 66.85 0.9225 ;
      LAYER metal3 ;
        RECT 66.78 0.055 66.85 1.4925 ;
      LAYER via1 ;
        RECT 66.7825 0.82 66.8475 0.885 ;
      LAYER via2 ;
        RECT 66.78 0.8175 66.85 0.8875 ;
    END
  END rs1_sel[9]
  PIN rs1_sel_bar[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 91.1525 0.9075 91.5025 0.9725 ;
        RECT 91.1525 0.8675 91.2225 1.0025 ;
      LAYER metal2 ;
        RECT 91.1525 0.865 91.2225 1.005 ;
      LAYER metal3 ;
        RECT 91.1525 0.055 91.2225 1.4925 ;
      LAYER via1 ;
        RECT 91.155 0.9025 91.22 0.9675 ;
      LAYER via2 ;
        RECT 91.1525 0.9 91.2225 0.97 ;
    END
  END rs1_sel_bar[0]
  PIN rs1_sel_bar[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.3775 0.9075 63.7275 0.9725 ;
        RECT 63.3775 0.8675 63.4475 1.0025 ;
      LAYER metal2 ;
        RECT 63.3775 0.865 63.4475 1.005 ;
      LAYER metal3 ;
        RECT 63.3775 0.055 63.4475 1.4925 ;
      LAYER via1 ;
        RECT 63.38 0.9025 63.445 0.9675 ;
      LAYER via2 ;
        RECT 63.3775 0.9 63.4475 0.97 ;
    END
  END rs1_sel_bar[10]
  PIN rs1_sel_bar[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 60.47 0.9075 60.82 0.9725 ;
        RECT 60.47 0.8675 60.54 1.0025 ;
      LAYER metal2 ;
        RECT 60.47 0.865 60.54 1.005 ;
      LAYER metal3 ;
        RECT 60.47 0.055 60.54 1.4925 ;
      LAYER via1 ;
        RECT 60.4725 0.9025 60.5375 0.9675 ;
      LAYER via2 ;
        RECT 60.47 0.9 60.54 0.97 ;
    END
  END rs1_sel_bar[11]
  PIN rs1_sel_bar[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 57.5625 0.9075 57.9125 0.9725 ;
        RECT 57.5625 0.8675 57.6325 1.0025 ;
      LAYER metal2 ;
        RECT 57.5625 0.865 57.6325 1.005 ;
      LAYER metal3 ;
        RECT 57.5625 0.055 57.6325 1.4925 ;
      LAYER via1 ;
        RECT 57.565 0.9025 57.63 0.9675 ;
      LAYER via2 ;
        RECT 57.5625 0.9 57.6325 0.97 ;
    END
  END rs1_sel_bar[12]
  PIN rs1_sel_bar[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 54.655 0.9075 55.005 0.9725 ;
        RECT 54.655 0.8675 54.725 1.0025 ;
      LAYER metal2 ;
        RECT 54.655 0.865 54.725 1.005 ;
      LAYER metal3 ;
        RECT 54.655 0.055 54.725 1.4925 ;
      LAYER via1 ;
        RECT 54.6575 0.9025 54.7225 0.9675 ;
      LAYER via2 ;
        RECT 54.655 0.9 54.725 0.97 ;
    END
  END rs1_sel_bar[13]
  PIN rs1_sel_bar[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 51.7475 0.9075 52.0975 0.9725 ;
        RECT 51.7475 0.8675 51.8175 1.0025 ;
      LAYER metal2 ;
        RECT 51.7475 0.865 51.8175 1.005 ;
      LAYER metal3 ;
        RECT 51.7475 0.055 51.8175 1.4925 ;
      LAYER via1 ;
        RECT 51.75 0.9025 51.815 0.9675 ;
      LAYER via2 ;
        RECT 51.7475 0.9 51.8175 0.97 ;
    END
  END rs1_sel_bar[14]
  PIN rs1_sel_bar[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 48.84 0.9075 49.19 0.9725 ;
        RECT 48.84 0.8675 48.91 1.0025 ;
      LAYER metal2 ;
        RECT 48.84 0.865 48.91 1.005 ;
      LAYER metal3 ;
        RECT 48.84 0.055 48.91 1.4925 ;
      LAYER via1 ;
        RECT 48.8425 0.9025 48.9075 0.9675 ;
      LAYER via2 ;
        RECT 48.84 0.9 48.91 0.97 ;
    END
  END rs1_sel_bar[15]
  PIN rs1_sel_bar[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 45.9325 0.9075 46.2825 0.9725 ;
        RECT 45.9325 0.8675 46.0025 1.0025 ;
      LAYER metal2 ;
        RECT 45.9325 0.865 46.0025 1.005 ;
      LAYER metal3 ;
        RECT 45.9325 0.055 46.0025 1.4925 ;
      LAYER via1 ;
        RECT 45.935 0.9025 46 0.9675 ;
      LAYER via2 ;
        RECT 45.9325 0.9 46.0025 0.97 ;
    END
  END rs1_sel_bar[16]
  PIN rs1_sel_bar[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 43.025 0.9075 43.375 0.9725 ;
        RECT 43.025 0.8675 43.095 1.0025 ;
      LAYER metal2 ;
        RECT 43.025 0.865 43.095 1.005 ;
      LAYER metal3 ;
        RECT 43.025 0.055 43.095 1.4925 ;
      LAYER via1 ;
        RECT 43.0275 0.9025 43.0925 0.9675 ;
      LAYER via2 ;
        RECT 43.025 0.9 43.095 0.97 ;
    END
  END rs1_sel_bar[17]
  PIN rs1_sel_bar[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 40.1175 0.9075 40.4675 0.9725 ;
        RECT 40.1175 0.8675 40.1875 1.0025 ;
      LAYER metal2 ;
        RECT 40.1175 0.865 40.1875 1.005 ;
      LAYER metal3 ;
        RECT 40.1175 0.055 40.1875 1.4925 ;
      LAYER via1 ;
        RECT 40.12 0.9025 40.185 0.9675 ;
      LAYER via2 ;
        RECT 40.1175 0.9 40.1875 0.97 ;
    END
  END rs1_sel_bar[18]
  PIN rs1_sel_bar[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 37.21 0.9075 37.56 0.9725 ;
        RECT 37.21 0.8675 37.28 1.0025 ;
      LAYER metal2 ;
        RECT 37.21 0.865 37.28 1.005 ;
      LAYER metal3 ;
        RECT 37.21 0.055 37.28 1.4925 ;
      LAYER via1 ;
        RECT 37.2125 0.9025 37.2775 0.9675 ;
      LAYER via2 ;
        RECT 37.21 0.9 37.28 0.97 ;
    END
  END rs1_sel_bar[19]
  PIN rs1_sel_bar[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 89.545 0.9075 89.895 0.9725 ;
        RECT 89.545 0.8675 89.615 1.0025 ;
      LAYER metal2 ;
        RECT 89.545 0.865 89.615 1.005 ;
      LAYER metal3 ;
        RECT 89.545 0.055 89.615 1.4925 ;
      LAYER via1 ;
        RECT 89.5475 0.9025 89.6125 0.9675 ;
      LAYER via2 ;
        RECT 89.545 0.9 89.615 0.97 ;
    END
  END rs1_sel_bar[1]
  PIN rs1_sel_bar[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 34.3025 0.9075 34.6525 0.9725 ;
        RECT 34.3025 0.8675 34.3725 1.0025 ;
      LAYER metal2 ;
        RECT 34.3025 0.865 34.3725 1.005 ;
      LAYER metal3 ;
        RECT 34.3025 0.055 34.3725 1.4925 ;
      LAYER via1 ;
        RECT 34.305 0.9025 34.37 0.9675 ;
      LAYER via2 ;
        RECT 34.3025 0.9 34.3725 0.97 ;
    END
  END rs1_sel_bar[20]
  PIN rs1_sel_bar[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 31.395 0.9075 31.745 0.9725 ;
        RECT 31.395 0.8675 31.465 1.0025 ;
      LAYER metal2 ;
        RECT 31.395 0.865 31.465 1.005 ;
      LAYER metal3 ;
        RECT 31.395 0.055 31.465 1.4925 ;
      LAYER via1 ;
        RECT 31.3975 0.9025 31.4625 0.9675 ;
      LAYER via2 ;
        RECT 31.395 0.9 31.465 0.97 ;
    END
  END rs1_sel_bar[21]
  PIN rs1_sel_bar[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 28.4875 0.9075 28.8375 0.9725 ;
        RECT 28.4875 0.8675 28.5575 1.0025 ;
      LAYER metal2 ;
        RECT 28.4875 0.865 28.5575 1.005 ;
      LAYER metal3 ;
        RECT 28.4875 0.055 28.5575 1.4925 ;
      LAYER via1 ;
        RECT 28.49 0.9025 28.555 0.9675 ;
      LAYER via2 ;
        RECT 28.4875 0.9 28.5575 0.97 ;
    END
  END rs1_sel_bar[22]
  PIN rs1_sel_bar[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 25.58 0.9075 25.93 0.9725 ;
        RECT 25.58 0.8675 25.65 1.0025 ;
      LAYER metal2 ;
        RECT 25.58 0.865 25.65 1.005 ;
      LAYER metal3 ;
        RECT 25.58 0.055 25.65 1.4925 ;
      LAYER via1 ;
        RECT 25.5825 0.9025 25.6475 0.9675 ;
      LAYER via2 ;
        RECT 25.58 0.9 25.65 0.97 ;
    END
  END rs1_sel_bar[23]
  PIN rs1_sel_bar[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 22.6725 0.9075 23.0225 0.9725 ;
        RECT 22.6725 0.8675 22.7425 1.0025 ;
      LAYER metal2 ;
        RECT 22.6725 0.865 22.7425 1.005 ;
      LAYER metal3 ;
        RECT 22.6725 0.055 22.7425 1.4925 ;
      LAYER via1 ;
        RECT 22.675 0.9025 22.74 0.9675 ;
      LAYER via2 ;
        RECT 22.6725 0.9 22.7425 0.97 ;
    END
  END rs1_sel_bar[24]
  PIN rs1_sel_bar[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 19.765 0.9075 20.115 0.9725 ;
        RECT 19.765 0.8675 19.835 1.0025 ;
      LAYER metal2 ;
        RECT 19.765 0.865 19.835 1.005 ;
      LAYER metal3 ;
        RECT 19.765 0.055 19.835 1.4925 ;
      LAYER via1 ;
        RECT 19.7675 0.9025 19.8325 0.9675 ;
      LAYER via2 ;
        RECT 19.765 0.9 19.835 0.97 ;
    END
  END rs1_sel_bar[25]
  PIN rs1_sel_bar[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 16.8575 0.9075 17.2075 0.9725 ;
        RECT 16.8575 0.8675 16.9275 1.0025 ;
      LAYER metal2 ;
        RECT 16.8575 0.865 16.9275 1.005 ;
      LAYER metal3 ;
        RECT 16.8575 0.055 16.9275 1.4925 ;
      LAYER via1 ;
        RECT 16.86 0.9025 16.925 0.9675 ;
      LAYER via2 ;
        RECT 16.8575 0.9 16.9275 0.97 ;
    END
  END rs1_sel_bar[26]
  PIN rs1_sel_bar[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 13.95 0.9075 14.3 0.9725 ;
        RECT 13.95 0.8675 14.02 1.0025 ;
      LAYER metal2 ;
        RECT 13.95 0.865 14.02 1.005 ;
      LAYER metal3 ;
        RECT 13.95 0.055 14.02 1.4925 ;
      LAYER via1 ;
        RECT 13.9525 0.9025 14.0175 0.9675 ;
      LAYER via2 ;
        RECT 13.95 0.9 14.02 0.97 ;
    END
  END rs1_sel_bar[27]
  PIN rs1_sel_bar[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 11.0425 0.9075 11.3925 0.9725 ;
        RECT 11.0425 0.8675 11.1125 1.0025 ;
      LAYER metal2 ;
        RECT 11.0425 0.865 11.1125 1.005 ;
      LAYER metal3 ;
        RECT 11.0425 0.055 11.1125 1.4925 ;
      LAYER via1 ;
        RECT 11.045 0.9025 11.11 0.9675 ;
      LAYER via2 ;
        RECT 11.0425 0.9 11.1125 0.97 ;
    END
  END rs1_sel_bar[28]
  PIN rs1_sel_bar[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 8.135 0.9075 8.485 0.9725 ;
        RECT 8.135 0.8675 8.205 1.0025 ;
      LAYER metal2 ;
        RECT 8.135 0.865 8.205 1.005 ;
      LAYER metal3 ;
        RECT 8.135 0.055 8.205 1.4925 ;
      LAYER via1 ;
        RECT 8.1375 0.9025 8.2025 0.9675 ;
      LAYER via2 ;
        RECT 8.135 0.9 8.205 0.97 ;
    END
  END rs1_sel_bar[29]
  PIN rs1_sel_bar[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 86.6375 0.9075 86.9875 0.9725 ;
        RECT 86.6375 0.8675 86.7075 1.0025 ;
      LAYER metal2 ;
        RECT 86.6375 0.865 86.7075 1.005 ;
      LAYER metal3 ;
        RECT 86.6375 0.055 86.7075 1.4925 ;
      LAYER via1 ;
        RECT 86.64 0.9025 86.705 0.9675 ;
      LAYER via2 ;
        RECT 86.6375 0.9 86.7075 0.97 ;
    END
  END rs1_sel_bar[2]
  PIN rs1_sel_bar[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.2275 0.9075 5.5775 0.9725 ;
        RECT 5.2275 0.8675 5.2975 1.0025 ;
      LAYER metal2 ;
        RECT 5.2275 0.865 5.2975 1.005 ;
      LAYER metal3 ;
        RECT 5.2275 0.055 5.2975 1.4925 ;
      LAYER via1 ;
        RECT 5.23 0.9025 5.295 0.9675 ;
      LAYER via2 ;
        RECT 5.2275 0.9 5.2975 0.97 ;
    END
  END rs1_sel_bar[30]
  PIN rs1_sel_bar[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.32 0.9075 2.67 0.9725 ;
        RECT 2.32 0.8675 2.39 1.0025 ;
      LAYER metal2 ;
        RECT 2.32 0.865 2.39 1.005 ;
      LAYER metal3 ;
        RECT 2.32 0.055 2.39 1.4925 ;
      LAYER via1 ;
        RECT 2.3225 0.9025 2.3875 0.9675 ;
      LAYER via2 ;
        RECT 2.32 0.9 2.39 0.97 ;
    END
  END rs1_sel_bar[31]
  PIN rs1_sel_bar[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 83.73 0.9075 84.08 0.9725 ;
        RECT 83.73 0.8675 83.8 1.0025 ;
      LAYER metal2 ;
        RECT 83.73 0.865 83.8 1.005 ;
      LAYER metal3 ;
        RECT 83.73 0.055 83.8 1.4925 ;
      LAYER via1 ;
        RECT 83.7325 0.9025 83.7975 0.9675 ;
      LAYER via2 ;
        RECT 83.73 0.9 83.8 0.97 ;
    END
  END rs1_sel_bar[3]
  PIN rs1_sel_bar[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 80.8225 0.9075 81.1725 0.9725 ;
        RECT 80.8225 0.8675 80.8925 1.0025 ;
      LAYER metal2 ;
        RECT 80.8225 0.865 80.8925 1.005 ;
      LAYER metal3 ;
        RECT 80.8225 0.055 80.8925 1.4925 ;
      LAYER via1 ;
        RECT 80.825 0.9025 80.89 0.9675 ;
      LAYER via2 ;
        RECT 80.8225 0.9 80.8925 0.97 ;
    END
  END rs1_sel_bar[4]
  PIN rs1_sel_bar[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 77.915 0.9075 78.265 0.9725 ;
        RECT 77.915 0.8675 77.985 1.0025 ;
      LAYER metal2 ;
        RECT 77.915 0.865 77.985 1.005 ;
      LAYER metal3 ;
        RECT 77.915 0.055 77.985 1.4925 ;
      LAYER via1 ;
        RECT 77.9175 0.9025 77.9825 0.9675 ;
      LAYER via2 ;
        RECT 77.915 0.9 77.985 0.97 ;
    END
  END rs1_sel_bar[5]
  PIN rs1_sel_bar[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 75.0075 0.9075 75.3575 0.9725 ;
        RECT 75.0075 0.8675 75.0775 1.0025 ;
      LAYER metal2 ;
        RECT 75.0075 0.865 75.0775 1.005 ;
      LAYER metal3 ;
        RECT 75.0075 0.055 75.0775 1.4925 ;
      LAYER via1 ;
        RECT 75.01 0.9025 75.075 0.9675 ;
      LAYER via2 ;
        RECT 75.0075 0.9 75.0775 0.97 ;
    END
  END rs1_sel_bar[6]
  PIN rs1_sel_bar[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 72.1 0.9075 72.45 0.9725 ;
        RECT 72.1 0.8675 72.17 1.0025 ;
      LAYER metal2 ;
        RECT 72.1 0.865 72.17 1.005 ;
      LAYER metal3 ;
        RECT 72.1 0.055 72.17 1.4925 ;
      LAYER via1 ;
        RECT 72.1025 0.9025 72.1675 0.9675 ;
      LAYER via2 ;
        RECT 72.1 0.9 72.17 0.97 ;
    END
  END rs1_sel_bar[7]
  PIN rs1_sel_bar[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 69.1925 0.9075 69.5425 0.9725 ;
        RECT 69.1925 0.8675 69.2625 1.0025 ;
      LAYER metal2 ;
        RECT 69.1925 0.865 69.2625 1.005 ;
      LAYER metal3 ;
        RECT 69.1925 0.055 69.2625 1.4925 ;
      LAYER via1 ;
        RECT 69.195 0.9025 69.26 0.9675 ;
      LAYER via2 ;
        RECT 69.1925 0.9 69.2625 0.97 ;
    END
  END rs1_sel_bar[8]
  PIN rs1_sel_bar[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 66.285 0.9075 66.635 0.9725 ;
        RECT 66.285 0.8675 66.355 1.0025 ;
      LAYER metal2 ;
        RECT 66.285 0.865 66.355 1.005 ;
      LAYER metal3 ;
        RECT 66.285 0.055 66.355 1.4925 ;
      LAYER via1 ;
        RECT 66.2875 0.9025 66.3525 0.9675 ;
      LAYER via2 ;
        RECT 66.285 0.9 66.355 0.97 ;
    END
  END rs1_sel_bar[9]
  PIN rs2_rdata
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 95.675 0.5825 95.745 0.7175 ;
        RECT 95.675 0.265 95.74 1.285 ;
        RECT 95.42 0.5325 95.74 0.5975 ;
        RECT 95.42 0.4975 95.485 0.6325 ;
      LAYER metal2 ;
        RECT 95.675 0.58 95.745 0.72 ;
      LAYER metal3 ;
        RECT 95.675 0.055 95.745 1.4925 ;
      LAYER via1 ;
        RECT 95.6775 0.6175 95.7425 0.6825 ;
      LAYER via2 ;
        RECT 95.675 0.615 95.745 0.685 ;
    END
  END rs2_rdata
  PIN rs2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 90.99 0.445 91.06 0.58 ;
        RECT 90.71 0.485 91.06 0.55 ;
      LAYER metal2 ;
        RECT 90.99 0.4425 91.06 0.5825 ;
      LAYER metal3 ;
        RECT 90.99 0.055 91.06 1.4925 ;
      LAYER via1 ;
        RECT 90.9925 0.48 91.0575 0.545 ;
      LAYER via2 ;
        RECT 90.99 0.4775 91.06 0.5475 ;
    END
  END rs2_sel[0]
  PIN rs2_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.215 0.445 63.285 0.58 ;
        RECT 62.935 0.485 63.285 0.55 ;
      LAYER metal2 ;
        RECT 63.215 0.4425 63.285 0.5825 ;
      LAYER metal3 ;
        RECT 63.215 0.055 63.285 1.4925 ;
      LAYER via1 ;
        RECT 63.2175 0.48 63.2825 0.545 ;
      LAYER via2 ;
        RECT 63.215 0.4775 63.285 0.5475 ;
    END
  END rs2_sel[10]
  PIN rs2_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 60.3075 0.445 60.3775 0.58 ;
        RECT 60.0275 0.485 60.3775 0.55 ;
      LAYER metal2 ;
        RECT 60.3075 0.4425 60.3775 0.5825 ;
      LAYER metal3 ;
        RECT 60.3075 0.055 60.3775 1.4925 ;
      LAYER via1 ;
        RECT 60.31 0.48 60.375 0.545 ;
      LAYER via2 ;
        RECT 60.3075 0.4775 60.3775 0.5475 ;
    END
  END rs2_sel[11]
  PIN rs2_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 57.4 0.445 57.47 0.58 ;
        RECT 57.12 0.485 57.47 0.55 ;
      LAYER metal2 ;
        RECT 57.4 0.4425 57.47 0.5825 ;
      LAYER metal3 ;
        RECT 57.4 0.055 57.47 1.4925 ;
      LAYER via1 ;
        RECT 57.4025 0.48 57.4675 0.545 ;
      LAYER via2 ;
        RECT 57.4 0.4775 57.47 0.5475 ;
    END
  END rs2_sel[12]
  PIN rs2_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 54.4925 0.445 54.5625 0.58 ;
        RECT 54.2125 0.485 54.5625 0.55 ;
      LAYER metal2 ;
        RECT 54.4925 0.4425 54.5625 0.5825 ;
      LAYER metal3 ;
        RECT 54.4925 0.055 54.5625 1.4925 ;
      LAYER via1 ;
        RECT 54.495 0.48 54.56 0.545 ;
      LAYER via2 ;
        RECT 54.4925 0.4775 54.5625 0.5475 ;
    END
  END rs2_sel[13]
  PIN rs2_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 51.585 0.445 51.655 0.58 ;
        RECT 51.305 0.485 51.655 0.55 ;
      LAYER metal2 ;
        RECT 51.585 0.4425 51.655 0.5825 ;
      LAYER metal3 ;
        RECT 51.585 0.055 51.655 1.4925 ;
      LAYER via1 ;
        RECT 51.5875 0.48 51.6525 0.545 ;
      LAYER via2 ;
        RECT 51.585 0.4775 51.655 0.5475 ;
    END
  END rs2_sel[14]
  PIN rs2_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 48.6775 0.445 48.7475 0.58 ;
        RECT 48.3975 0.485 48.7475 0.55 ;
      LAYER metal2 ;
        RECT 48.6775 0.4425 48.7475 0.5825 ;
      LAYER metal3 ;
        RECT 48.6775 0.055 48.7475 1.4925 ;
      LAYER via1 ;
        RECT 48.68 0.48 48.745 0.545 ;
      LAYER via2 ;
        RECT 48.6775 0.4775 48.7475 0.5475 ;
    END
  END rs2_sel[15]
  PIN rs2_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 45.77 0.445 45.84 0.58 ;
        RECT 45.49 0.485 45.84 0.55 ;
      LAYER metal2 ;
        RECT 45.77 0.4425 45.84 0.5825 ;
      LAYER metal3 ;
        RECT 45.77 0.055 45.84 1.4925 ;
      LAYER via1 ;
        RECT 45.7725 0.48 45.8375 0.545 ;
      LAYER via2 ;
        RECT 45.77 0.4775 45.84 0.5475 ;
    END
  END rs2_sel[16]
  PIN rs2_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 42.8625 0.445 42.9325 0.58 ;
        RECT 42.5825 0.485 42.9325 0.55 ;
      LAYER metal2 ;
        RECT 42.8625 0.4425 42.9325 0.5825 ;
      LAYER metal3 ;
        RECT 42.8625 0.055 42.9325 1.4925 ;
      LAYER via1 ;
        RECT 42.865 0.48 42.93 0.545 ;
      LAYER via2 ;
        RECT 42.8625 0.4775 42.9325 0.5475 ;
    END
  END rs2_sel[17]
  PIN rs2_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 39.955 0.445 40.025 0.58 ;
        RECT 39.675 0.485 40.025 0.55 ;
      LAYER metal2 ;
        RECT 39.955 0.4425 40.025 0.5825 ;
      LAYER metal3 ;
        RECT 39.955 0.055 40.025 1.4925 ;
      LAYER via1 ;
        RECT 39.9575 0.48 40.0225 0.545 ;
      LAYER via2 ;
        RECT 39.955 0.4775 40.025 0.5475 ;
    END
  END rs2_sel[18]
  PIN rs2_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 37.0475 0.445 37.1175 0.58 ;
        RECT 36.7675 0.485 37.1175 0.55 ;
      LAYER metal2 ;
        RECT 37.0475 0.4425 37.1175 0.5825 ;
      LAYER metal3 ;
        RECT 37.0475 0.055 37.1175 1.4925 ;
      LAYER via1 ;
        RECT 37.05 0.48 37.115 0.545 ;
      LAYER via2 ;
        RECT 37.0475 0.4775 37.1175 0.5475 ;
    END
  END rs2_sel[19]
  PIN rs2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 89.3825 0.445 89.4525 0.58 ;
        RECT 89.1025 0.485 89.4525 0.55 ;
      LAYER metal2 ;
        RECT 89.3825 0.4425 89.4525 0.5825 ;
      LAYER metal3 ;
        RECT 89.3825 0.055 89.4525 1.4925 ;
      LAYER via1 ;
        RECT 89.385 0.48 89.45 0.545 ;
      LAYER via2 ;
        RECT 89.3825 0.4775 89.4525 0.5475 ;
    END
  END rs2_sel[1]
  PIN rs2_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 34.14 0.445 34.21 0.58 ;
        RECT 33.86 0.485 34.21 0.55 ;
      LAYER metal2 ;
        RECT 34.14 0.4425 34.21 0.5825 ;
      LAYER metal3 ;
        RECT 34.14 0.055 34.21 1.4925 ;
      LAYER via1 ;
        RECT 34.1425 0.48 34.2075 0.545 ;
      LAYER via2 ;
        RECT 34.14 0.4775 34.21 0.5475 ;
    END
  END rs2_sel[20]
  PIN rs2_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 31.2325 0.445 31.3025 0.58 ;
        RECT 30.9525 0.485 31.3025 0.55 ;
      LAYER metal2 ;
        RECT 31.2325 0.4425 31.3025 0.5825 ;
      LAYER metal3 ;
        RECT 31.2325 0.055 31.3025 1.4925 ;
      LAYER via1 ;
        RECT 31.235 0.48 31.3 0.545 ;
      LAYER via2 ;
        RECT 31.2325 0.4775 31.3025 0.5475 ;
    END
  END rs2_sel[21]
  PIN rs2_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 28.325 0.445 28.395 0.58 ;
        RECT 28.045 0.485 28.395 0.55 ;
      LAYER metal2 ;
        RECT 28.325 0.4425 28.395 0.5825 ;
      LAYER metal3 ;
        RECT 28.325 0.055 28.395 1.4925 ;
      LAYER via1 ;
        RECT 28.3275 0.48 28.3925 0.545 ;
      LAYER via2 ;
        RECT 28.325 0.4775 28.395 0.5475 ;
    END
  END rs2_sel[22]
  PIN rs2_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 25.4175 0.445 25.4875 0.58 ;
        RECT 25.1375 0.485 25.4875 0.55 ;
      LAYER metal2 ;
        RECT 25.4175 0.4425 25.4875 0.5825 ;
      LAYER metal3 ;
        RECT 25.4175 0.055 25.4875 1.4925 ;
      LAYER via1 ;
        RECT 25.42 0.48 25.485 0.545 ;
      LAYER via2 ;
        RECT 25.4175 0.4775 25.4875 0.5475 ;
    END
  END rs2_sel[23]
  PIN rs2_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 22.51 0.445 22.58 0.58 ;
        RECT 22.23 0.485 22.58 0.55 ;
      LAYER metal2 ;
        RECT 22.51 0.4425 22.58 0.5825 ;
      LAYER metal3 ;
        RECT 22.51 0.055 22.58 1.4925 ;
      LAYER via1 ;
        RECT 22.5125 0.48 22.5775 0.545 ;
      LAYER via2 ;
        RECT 22.51 0.4775 22.58 0.5475 ;
    END
  END rs2_sel[24]
  PIN rs2_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 19.6025 0.445 19.6725 0.58 ;
        RECT 19.3225 0.485 19.6725 0.55 ;
      LAYER metal2 ;
        RECT 19.6025 0.4425 19.6725 0.5825 ;
      LAYER metal3 ;
        RECT 19.6025 0.055 19.6725 1.4925 ;
      LAYER via1 ;
        RECT 19.605 0.48 19.67 0.545 ;
      LAYER via2 ;
        RECT 19.6025 0.4775 19.6725 0.5475 ;
    END
  END rs2_sel[25]
  PIN rs2_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 16.695 0.445 16.765 0.58 ;
        RECT 16.415 0.485 16.765 0.55 ;
      LAYER metal2 ;
        RECT 16.695 0.4425 16.765 0.5825 ;
      LAYER metal3 ;
        RECT 16.695 0.055 16.765 1.4925 ;
      LAYER via1 ;
        RECT 16.6975 0.48 16.7625 0.545 ;
      LAYER via2 ;
        RECT 16.695 0.4775 16.765 0.5475 ;
    END
  END rs2_sel[26]
  PIN rs2_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 13.7875 0.445 13.8575 0.58 ;
        RECT 13.5075 0.485 13.8575 0.55 ;
      LAYER metal2 ;
        RECT 13.7875 0.4425 13.8575 0.5825 ;
      LAYER metal3 ;
        RECT 13.7875 0.055 13.8575 1.4925 ;
      LAYER via1 ;
        RECT 13.79 0.48 13.855 0.545 ;
      LAYER via2 ;
        RECT 13.7875 0.4775 13.8575 0.5475 ;
    END
  END rs2_sel[27]
  PIN rs2_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 10.88 0.445 10.95 0.58 ;
        RECT 10.6 0.485 10.95 0.55 ;
      LAYER metal2 ;
        RECT 10.88 0.4425 10.95 0.5825 ;
      LAYER metal3 ;
        RECT 10.88 0.055 10.95 1.4925 ;
      LAYER via1 ;
        RECT 10.8825 0.48 10.9475 0.545 ;
      LAYER via2 ;
        RECT 10.88 0.4775 10.95 0.5475 ;
    END
  END rs2_sel[28]
  PIN rs2_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 7.9725 0.445 8.0425 0.58 ;
        RECT 7.6925 0.485 8.0425 0.55 ;
      LAYER metal2 ;
        RECT 7.9725 0.4425 8.0425 0.5825 ;
      LAYER metal3 ;
        RECT 7.9725 0.055 8.0425 1.4925 ;
      LAYER via1 ;
        RECT 7.975 0.48 8.04 0.545 ;
      LAYER via2 ;
        RECT 7.9725 0.4775 8.0425 0.5475 ;
    END
  END rs2_sel[29]
  PIN rs2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 86.475 0.445 86.545 0.58 ;
        RECT 86.195 0.485 86.545 0.55 ;
      LAYER metal2 ;
        RECT 86.475 0.4425 86.545 0.5825 ;
      LAYER metal3 ;
        RECT 86.475 0.055 86.545 1.4925 ;
      LAYER via1 ;
        RECT 86.4775 0.48 86.5425 0.545 ;
      LAYER via2 ;
        RECT 86.475 0.4775 86.545 0.5475 ;
    END
  END rs2_sel[2]
  PIN rs2_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.065 0.445 5.135 0.58 ;
        RECT 4.785 0.485 5.135 0.55 ;
      LAYER metal2 ;
        RECT 5.065 0.4425 5.135 0.5825 ;
      LAYER metal3 ;
        RECT 5.065 0.055 5.135 1.4925 ;
      LAYER via1 ;
        RECT 5.0675 0.48 5.1325 0.545 ;
      LAYER via2 ;
        RECT 5.065 0.4775 5.135 0.5475 ;
    END
  END rs2_sel[30]
  PIN rs2_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.1575 0.445 2.2275 0.58 ;
        RECT 1.8775 0.485 2.2275 0.55 ;
      LAYER metal2 ;
        RECT 2.1575 0.4425 2.2275 0.5825 ;
      LAYER metal3 ;
        RECT 2.1575 0.055 2.2275 1.49 ;
      LAYER via1 ;
        RECT 2.16 0.48 2.225 0.545 ;
      LAYER via2 ;
        RECT 2.1575 0.4775 2.2275 0.5475 ;
    END
  END rs2_sel[31]
  PIN rs2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 83.5675 0.445 83.6375 0.58 ;
        RECT 83.2875 0.485 83.6375 0.55 ;
      LAYER metal2 ;
        RECT 83.5675 0.4425 83.6375 0.5825 ;
      LAYER metal3 ;
        RECT 83.5675 0.055 83.6375 1.4925 ;
      LAYER via1 ;
        RECT 83.57 0.48 83.635 0.545 ;
      LAYER via2 ;
        RECT 83.5675 0.4775 83.6375 0.5475 ;
    END
  END rs2_sel[3]
  PIN rs2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 80.66 0.445 80.73 0.58 ;
        RECT 80.38 0.485 80.73 0.55 ;
      LAYER metal2 ;
        RECT 80.66 0.4425 80.73 0.5825 ;
      LAYER metal3 ;
        RECT 80.66 0.055 80.73 1.4925 ;
      LAYER via1 ;
        RECT 80.6625 0.48 80.7275 0.545 ;
      LAYER via2 ;
        RECT 80.66 0.4775 80.73 0.5475 ;
    END
  END rs2_sel[4]
  PIN rs2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 77.7525 0.445 77.8225 0.58 ;
        RECT 77.4725 0.485 77.8225 0.55 ;
      LAYER metal2 ;
        RECT 77.7525 0.4425 77.8225 0.5825 ;
      LAYER metal3 ;
        RECT 77.7525 0.055 77.8225 1.4925 ;
      LAYER via1 ;
        RECT 77.755 0.48 77.82 0.545 ;
      LAYER via2 ;
        RECT 77.7525 0.4775 77.8225 0.5475 ;
    END
  END rs2_sel[5]
  PIN rs2_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 74.845 0.445 74.915 0.58 ;
        RECT 74.565 0.485 74.915 0.55 ;
      LAYER metal2 ;
        RECT 74.845 0.4425 74.915 0.5825 ;
      LAYER metal3 ;
        RECT 74.845 0.055 74.915 1.4925 ;
      LAYER via1 ;
        RECT 74.8475 0.48 74.9125 0.545 ;
      LAYER via2 ;
        RECT 74.845 0.4775 74.915 0.5475 ;
    END
  END rs2_sel[6]
  PIN rs2_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 71.9375 0.445 72.0075 0.58 ;
        RECT 71.6575 0.485 72.0075 0.55 ;
      LAYER metal2 ;
        RECT 71.9375 0.4425 72.0075 0.5825 ;
      LAYER metal3 ;
        RECT 71.9375 0.055 72.0075 1.4925 ;
      LAYER via1 ;
        RECT 71.94 0.48 72.005 0.545 ;
      LAYER via2 ;
        RECT 71.9375 0.4775 72.0075 0.5475 ;
    END
  END rs2_sel[7]
  PIN rs2_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 69.03 0.445 69.1 0.58 ;
        RECT 68.75 0.485 69.1 0.55 ;
      LAYER metal2 ;
        RECT 69.03 0.4425 69.1 0.5825 ;
      LAYER metal3 ;
        RECT 69.03 0.055 69.1 1.4925 ;
      LAYER via1 ;
        RECT 69.0325 0.48 69.0975 0.545 ;
      LAYER via2 ;
        RECT 69.03 0.4775 69.1 0.5475 ;
    END
  END rs2_sel[8]
  PIN rs2_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 66.1225 0.445 66.1925 0.58 ;
        RECT 65.8425 0.485 66.1925 0.55 ;
      LAYER metal2 ;
        RECT 66.1225 0.4425 66.1925 0.5825 ;
      LAYER metal3 ;
        RECT 66.1225 0.055 66.1925 1.4925 ;
      LAYER via1 ;
        RECT 66.125 0.48 66.19 0.545 ;
      LAYER via2 ;
        RECT 66.1225 0.4775 66.1925 0.5475 ;
    END
  END rs2_sel[9]
  PIN rs2_sel_bar[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 90.5075 0.9075 90.845 0.9725 ;
        RECT 90.5075 0.8675 90.5775 1.0025 ;
      LAYER metal2 ;
        RECT 90.5075 0.865 90.5775 1.005 ;
      LAYER metal3 ;
        RECT 90.5075 0.055 90.5775 1.4925 ;
      LAYER via1 ;
        RECT 90.51 0.9025 90.575 0.9675 ;
      LAYER via2 ;
        RECT 90.5075 0.9 90.5775 0.97 ;
    END
  END rs2_sel_bar[0]
  PIN rs2_sel_bar[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 62.7325 0.9075 63.07 0.9725 ;
        RECT 62.7325 0.8675 62.8025 1.0025 ;
      LAYER metal2 ;
        RECT 62.7325 0.865 62.8025 1.005 ;
      LAYER metal3 ;
        RECT 62.7325 0.055 62.8025 1.4925 ;
      LAYER via1 ;
        RECT 62.735 0.9025 62.8 0.9675 ;
      LAYER via2 ;
        RECT 62.7325 0.9 62.8025 0.97 ;
    END
  END rs2_sel_bar[10]
  PIN rs2_sel_bar[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 59.825 0.9075 60.1625 0.9725 ;
        RECT 59.825 0.8675 59.895 1.0025 ;
      LAYER metal2 ;
        RECT 59.825 0.865 59.895 1.005 ;
      LAYER metal3 ;
        RECT 59.825 0.055 59.895 1.4925 ;
      LAYER via1 ;
        RECT 59.8275 0.9025 59.8925 0.9675 ;
      LAYER via2 ;
        RECT 59.825 0.9 59.895 0.97 ;
    END
  END rs2_sel_bar[11]
  PIN rs2_sel_bar[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 56.9175 0.9075 57.255 0.9725 ;
        RECT 56.9175 0.8675 56.9875 1.0025 ;
      LAYER metal2 ;
        RECT 56.9175 0.865 56.9875 1.005 ;
      LAYER metal3 ;
        RECT 56.9175 0.055 56.9875 1.4925 ;
      LAYER via1 ;
        RECT 56.92 0.9025 56.985 0.9675 ;
      LAYER via2 ;
        RECT 56.9175 0.9 56.9875 0.97 ;
    END
  END rs2_sel_bar[12]
  PIN rs2_sel_bar[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 54.01 0.9075 54.3475 0.9725 ;
        RECT 54.01 0.8675 54.08 1.0025 ;
      LAYER metal2 ;
        RECT 54.01 0.865 54.08 1.005 ;
      LAYER metal3 ;
        RECT 54.01 0.055 54.08 1.4925 ;
      LAYER via1 ;
        RECT 54.0125 0.9025 54.0775 0.9675 ;
      LAYER via2 ;
        RECT 54.01 0.9 54.08 0.97 ;
    END
  END rs2_sel_bar[13]
  PIN rs2_sel_bar[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 51.1025 0.9075 51.44 0.9725 ;
        RECT 51.1025 0.8675 51.1725 1.0025 ;
      LAYER metal2 ;
        RECT 51.1025 0.865 51.1725 1.005 ;
      LAYER metal3 ;
        RECT 51.1025 0.055 51.1725 1.4925 ;
      LAYER via1 ;
        RECT 51.105 0.9025 51.17 0.9675 ;
      LAYER via2 ;
        RECT 51.1025 0.9 51.1725 0.97 ;
    END
  END rs2_sel_bar[14]
  PIN rs2_sel_bar[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 48.195 0.9075 48.5325 0.9725 ;
        RECT 48.195 0.8675 48.265 1.0025 ;
      LAYER metal2 ;
        RECT 48.195 0.865 48.265 1.005 ;
      LAYER metal3 ;
        RECT 48.195 0.055 48.265 1.4925 ;
      LAYER via1 ;
        RECT 48.1975 0.9025 48.2625 0.9675 ;
      LAYER via2 ;
        RECT 48.195 0.9 48.265 0.97 ;
    END
  END rs2_sel_bar[15]
  PIN rs2_sel_bar[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 45.2875 0.9075 45.625 0.9725 ;
        RECT 45.2875 0.8675 45.3575 1.0025 ;
      LAYER metal2 ;
        RECT 45.2875 0.865 45.3575 1.005 ;
      LAYER metal3 ;
        RECT 45.2875 0.055 45.3575 1.4925 ;
      LAYER via1 ;
        RECT 45.29 0.9025 45.355 0.9675 ;
      LAYER via2 ;
        RECT 45.2875 0.9 45.3575 0.97 ;
    END
  END rs2_sel_bar[16]
  PIN rs2_sel_bar[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 42.38 0.9075 42.7175 0.9725 ;
        RECT 42.38 0.8675 42.45 1.0025 ;
      LAYER metal2 ;
        RECT 42.38 0.865 42.45 1.005 ;
      LAYER metal3 ;
        RECT 42.38 0.055 42.45 1.4925 ;
      LAYER via1 ;
        RECT 42.3825 0.9025 42.4475 0.9675 ;
      LAYER via2 ;
        RECT 42.38 0.9 42.45 0.97 ;
    END
  END rs2_sel_bar[17]
  PIN rs2_sel_bar[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 39.4725 0.9075 39.81 0.9725 ;
        RECT 39.4725 0.8675 39.5425 1.0025 ;
      LAYER metal2 ;
        RECT 39.4725 0.865 39.5425 1.005 ;
      LAYER metal3 ;
        RECT 39.4725 0.055 39.5425 1.4925 ;
      LAYER via1 ;
        RECT 39.475 0.9025 39.54 0.9675 ;
      LAYER via2 ;
        RECT 39.4725 0.9 39.5425 0.97 ;
    END
  END rs2_sel_bar[18]
  PIN rs2_sel_bar[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 36.565 0.9075 36.9025 0.9725 ;
        RECT 36.565 0.8675 36.635 1.0025 ;
      LAYER metal2 ;
        RECT 36.565 0.865 36.635 1.005 ;
      LAYER metal3 ;
        RECT 36.565 0.055 36.635 1.4925 ;
      LAYER via1 ;
        RECT 36.5675 0.9025 36.6325 0.9675 ;
      LAYER via2 ;
        RECT 36.565 0.9 36.635 0.97 ;
    END
  END rs2_sel_bar[19]
  PIN rs2_sel_bar[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 88.9 0.9075 89.2375 0.9725 ;
        RECT 88.9 0.8675 88.97 1.0025 ;
      LAYER metal2 ;
        RECT 88.9 0.865 88.97 1.005 ;
      LAYER metal3 ;
        RECT 88.9 0.055 88.97 1.4925 ;
      LAYER via1 ;
        RECT 88.9025 0.9025 88.9675 0.9675 ;
      LAYER via2 ;
        RECT 88.9 0.9 88.97 0.97 ;
    END
  END rs2_sel_bar[1]
  PIN rs2_sel_bar[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 33.6575 0.9075 33.995 0.9725 ;
        RECT 33.6575 0.8675 33.7275 1.0025 ;
      LAYER metal2 ;
        RECT 33.6575 0.865 33.7275 1.005 ;
      LAYER metal3 ;
        RECT 33.6575 0.055 33.7275 1.4925 ;
      LAYER via1 ;
        RECT 33.66 0.9025 33.725 0.9675 ;
      LAYER via2 ;
        RECT 33.6575 0.9 33.7275 0.97 ;
    END
  END rs2_sel_bar[20]
  PIN rs2_sel_bar[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 30.75 0.9075 31.0875 0.9725 ;
        RECT 30.75 0.8675 30.82 1.0025 ;
      LAYER metal2 ;
        RECT 30.75 0.865 30.82 1.005 ;
      LAYER metal3 ;
        RECT 30.75 0.055 30.82 1.4925 ;
      LAYER via1 ;
        RECT 30.7525 0.9025 30.8175 0.9675 ;
      LAYER via2 ;
        RECT 30.75 0.9 30.82 0.97 ;
    END
  END rs2_sel_bar[21]
  PIN rs2_sel_bar[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 27.8425 0.9075 28.18 0.9725 ;
        RECT 27.8425 0.8675 27.9125 1.0025 ;
      LAYER metal2 ;
        RECT 27.8425 0.865 27.9125 1.005 ;
      LAYER metal3 ;
        RECT 27.8425 0.055 27.9125 1.4925 ;
      LAYER via1 ;
        RECT 27.845 0.9025 27.91 0.9675 ;
      LAYER via2 ;
        RECT 27.8425 0.9 27.9125 0.97 ;
    END
  END rs2_sel_bar[22]
  PIN rs2_sel_bar[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 24.935 0.9075 25.2725 0.9725 ;
        RECT 24.935 0.8675 25.005 1.0025 ;
      LAYER metal2 ;
        RECT 24.935 0.865 25.005 1.005 ;
      LAYER metal3 ;
        RECT 24.935 0.055 25.005 1.4925 ;
      LAYER via1 ;
        RECT 24.9375 0.9025 25.0025 0.9675 ;
      LAYER via2 ;
        RECT 24.935 0.9 25.005 0.97 ;
    END
  END rs2_sel_bar[23]
  PIN rs2_sel_bar[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 22.0275 0.9075 22.365 0.9725 ;
        RECT 22.0275 0.8675 22.0975 1.0025 ;
      LAYER metal2 ;
        RECT 22.0275 0.865 22.0975 1.005 ;
      LAYER metal3 ;
        RECT 22.0275 0.055 22.0975 1.4925 ;
      LAYER via1 ;
        RECT 22.03 0.9025 22.095 0.9675 ;
      LAYER via2 ;
        RECT 22.0275 0.9 22.0975 0.97 ;
    END
  END rs2_sel_bar[24]
  PIN rs2_sel_bar[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 19.12 0.9075 19.4575 0.9725 ;
        RECT 19.12 0.8675 19.19 1.0025 ;
      LAYER metal2 ;
        RECT 19.12 0.865 19.19 1.005 ;
      LAYER metal3 ;
        RECT 19.12 0.055 19.19 1.4925 ;
      LAYER via1 ;
        RECT 19.1225 0.9025 19.1875 0.9675 ;
      LAYER via2 ;
        RECT 19.12 0.9 19.19 0.97 ;
    END
  END rs2_sel_bar[25]
  PIN rs2_sel_bar[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 16.2125 0.9075 16.55 0.9725 ;
        RECT 16.2125 0.8675 16.2825 1.0025 ;
      LAYER metal2 ;
        RECT 16.2125 0.865 16.2825 1.005 ;
      LAYER metal3 ;
        RECT 16.2125 0.055 16.2825 1.4925 ;
      LAYER via1 ;
        RECT 16.215 0.9025 16.28 0.9675 ;
      LAYER via2 ;
        RECT 16.2125 0.9 16.2825 0.97 ;
    END
  END rs2_sel_bar[26]
  PIN rs2_sel_bar[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 13.305 0.9075 13.6425 0.9725 ;
        RECT 13.305 0.8675 13.375 1.0025 ;
      LAYER metal2 ;
        RECT 13.305 0.865 13.375 1.005 ;
      LAYER metal3 ;
        RECT 13.305 0.055 13.375 1.4925 ;
      LAYER via1 ;
        RECT 13.3075 0.9025 13.3725 0.9675 ;
      LAYER via2 ;
        RECT 13.305 0.9 13.375 0.97 ;
    END
  END rs2_sel_bar[27]
  PIN rs2_sel_bar[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 10.3975 0.9075 10.735 0.9725 ;
        RECT 10.3975 0.8675 10.4675 1.0025 ;
      LAYER metal2 ;
        RECT 10.3975 0.865 10.4675 1.005 ;
      LAYER metal3 ;
        RECT 10.3975 0.055 10.4675 1.4925 ;
      LAYER via1 ;
        RECT 10.4 0.9025 10.465 0.9675 ;
      LAYER via2 ;
        RECT 10.3975 0.9 10.4675 0.97 ;
    END
  END rs2_sel_bar[28]
  PIN rs2_sel_bar[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 7.49 0.9075 7.8275 0.9725 ;
        RECT 7.49 0.8675 7.56 1.0025 ;
      LAYER metal2 ;
        RECT 7.49 0.865 7.56 1.005 ;
      LAYER metal3 ;
        RECT 7.49 0.055 7.56 1.4925 ;
      LAYER via1 ;
        RECT 7.4925 0.9025 7.5575 0.9675 ;
      LAYER via2 ;
        RECT 7.49 0.9 7.56 0.97 ;
    END
  END rs2_sel_bar[29]
  PIN rs2_sel_bar[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 85.9925 0.9075 86.33 0.9725 ;
        RECT 85.9925 0.8675 86.0625 1.0025 ;
      LAYER metal2 ;
        RECT 85.9925 0.865 86.0625 1.005 ;
      LAYER metal3 ;
        RECT 85.9925 0.055 86.0625 1.4925 ;
      LAYER via1 ;
        RECT 85.995 0.9025 86.06 0.9675 ;
      LAYER via2 ;
        RECT 85.9925 0.9 86.0625 0.97 ;
    END
  END rs2_sel_bar[2]
  PIN rs2_sel_bar[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.5825 0.9075 4.92 0.9725 ;
        RECT 4.5825 0.8675 4.6525 1.0025 ;
      LAYER metal2 ;
        RECT 4.5825 0.865 4.6525 1.005 ;
      LAYER metal3 ;
        RECT 4.5825 0.055 4.6525 1.4925 ;
      LAYER via1 ;
        RECT 4.585 0.9025 4.65 0.9675 ;
      LAYER via2 ;
        RECT 4.5825 0.9 4.6525 0.97 ;
    END
  END rs2_sel_bar[30]
  PIN rs2_sel_bar[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.675 0.9075 2.0125 0.9725 ;
        RECT 1.675 0.8675 1.745 1.0025 ;
      LAYER metal2 ;
        RECT 1.675 0.865 1.745 1.005 ;
      LAYER metal3 ;
        RECT 1.675 0.055 1.745 1.4925 ;
      LAYER via1 ;
        RECT 1.6775 0.9025 1.7425 0.9675 ;
      LAYER via2 ;
        RECT 1.675 0.9 1.745 0.97 ;
    END
  END rs2_sel_bar[31]
  PIN rs2_sel_bar[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 83.085 0.9075 83.4225 0.9725 ;
        RECT 83.085 0.8675 83.155 1.0025 ;
      LAYER metal2 ;
        RECT 83.085 0.865 83.155 1.005 ;
      LAYER metal3 ;
        RECT 83.085 0.055 83.155 1.4925 ;
      LAYER via1 ;
        RECT 83.0875 0.9025 83.1525 0.9675 ;
      LAYER via2 ;
        RECT 83.085 0.9 83.155 0.97 ;
    END
  END rs2_sel_bar[3]
  PIN rs2_sel_bar[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 80.1775 0.9075 80.515 0.9725 ;
        RECT 80.1775 0.8675 80.2475 1.0025 ;
      LAYER metal2 ;
        RECT 80.1775 0.865 80.2475 1.005 ;
      LAYER metal3 ;
        RECT 80.1775 0.055 80.2475 1.4925 ;
      LAYER via1 ;
        RECT 80.18 0.9025 80.245 0.9675 ;
      LAYER via2 ;
        RECT 80.1775 0.9 80.2475 0.97 ;
    END
  END rs2_sel_bar[4]
  PIN rs2_sel_bar[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 77.27 0.9075 77.6075 0.9725 ;
        RECT 77.27 0.8675 77.34 1.0025 ;
      LAYER metal2 ;
        RECT 77.27 0.865 77.34 1.005 ;
      LAYER metal3 ;
        RECT 77.27 0.055 77.34 1.4925 ;
      LAYER via1 ;
        RECT 77.2725 0.9025 77.3375 0.9675 ;
      LAYER via2 ;
        RECT 77.27 0.9 77.34 0.97 ;
    END
  END rs2_sel_bar[5]
  PIN rs2_sel_bar[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 74.3625 0.9075 74.7 0.9725 ;
        RECT 74.3625 0.8675 74.4325 1.0025 ;
      LAYER metal2 ;
        RECT 74.3625 0.865 74.4325 1.005 ;
      LAYER metal3 ;
        RECT 74.3625 0.055 74.4325 1.4925 ;
      LAYER via1 ;
        RECT 74.365 0.9025 74.43 0.9675 ;
      LAYER via2 ;
        RECT 74.3625 0.9 74.4325 0.97 ;
    END
  END rs2_sel_bar[6]
  PIN rs2_sel_bar[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 71.455 0.9075 71.7925 0.9725 ;
        RECT 71.455 0.8675 71.525 1.0025 ;
      LAYER metal2 ;
        RECT 71.455 0.865 71.525 1.005 ;
      LAYER metal3 ;
        RECT 71.455 0.055 71.525 1.4925 ;
      LAYER via1 ;
        RECT 71.4575 0.9025 71.5225 0.9675 ;
      LAYER via2 ;
        RECT 71.455 0.9 71.525 0.97 ;
    END
  END rs2_sel_bar[7]
  PIN rs2_sel_bar[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 68.5475 0.9075 68.885 0.9725 ;
        RECT 68.5475 0.8675 68.6175 1.0025 ;
      LAYER metal2 ;
        RECT 68.5475 0.865 68.6175 1.005 ;
      LAYER metal3 ;
        RECT 68.5475 0.055 68.6175 1.4925 ;
      LAYER via1 ;
        RECT 68.55 0.9025 68.615 0.9675 ;
      LAYER via2 ;
        RECT 68.5475 0.9 68.6175 0.97 ;
    END
  END rs2_sel_bar[8]
  PIN rs2_sel_bar[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 65.64 0.9075 65.9775 0.9725 ;
        RECT 65.64 0.8675 65.71 1.0025 ;
      LAYER metal2 ;
        RECT 65.64 0.865 65.71 1.005 ;
      LAYER metal3 ;
        RECT 65.64 0.055 65.71 1.4925 ;
      LAYER via1 ;
        RECT 65.6425 0.9025 65.7075 0.9675 ;
      LAYER via2 ;
        RECT 65.64 0.9 65.71 0.97 ;
    END
  END rs2_sel_bar[9]
  OBS
    LAYER metal1 ;
      RECT 95.0125 0.715 95.0775 0.85 ;
      RECT 95.0125 0.75 95.2625 0.815 ;
      RECT 95.1975 0.5125 95.2625 0.815 ;
      RECT 94.575 0.265 94.64 1.285 ;
      RECT 95.1975 0.88 95.2625 1.015 ;
      RECT 94.8775 0.915 95.2625 0.98 ;
      RECT 94.8775 0.55 94.9425 0.98 ;
      RECT 95.0125 0.515 95.0775 0.65 ;
      RECT 94.575 0.5525 94.9425 0.6175 ;
      RECT 94.8775 0.55 95.0775 0.615 ;
      RECT 94.2 0.265 94.265 1.285 ;
      RECT 94.4325 0.505 94.4975 0.64 ;
      RECT 94.2 0.54 94.4975 0.605 ;
      RECT 94.015 0.265 94.08 1.285 ;
      RECT 94.015 0.49 94.0825 0.625 ;
      RECT 92.9825 0.715 93.0475 0.85 ;
      RECT 92.9825 0.75 93.2325 0.815 ;
      RECT 93.1675 0.5125 93.2325 0.815 ;
      RECT 92.545 0.265 92.61 1.285 ;
      RECT 93.1675 0.88 93.2325 1.015 ;
      RECT 92.8475 0.915 93.2325 0.98 ;
      RECT 92.8475 0.55 92.9125 0.98 ;
      RECT 92.9825 0.515 93.0475 0.65 ;
      RECT 92.545 0.5525 92.9125 0.6175 ;
      RECT 92.8475 0.55 93.0475 0.615 ;
      RECT 92.17 0.265 92.235 1.285 ;
      RECT 92.4025 0.505 92.4675 0.64 ;
      RECT 92.17 0.54 92.4675 0.605 ;
      RECT 91.985 0.265 92.05 1.285 ;
      RECT 91.985 0.49 92.0525 0.625 ;
      RECT 91.495 1.0425 91.56 1.2825 ;
      RECT 91.4925 1.095 91.5625 1.235 ;
      RECT 90.3775 0.265 90.4425 1.285 ;
      RECT 91.31 0.6575 91.375 0.7925 ;
      RECT 90.6525 0.6475 90.7175 0.7825 ;
      RECT 90.6525 0.685 91.375 0.75 ;
      RECT 90.3775 0.6825 90.7175 0.7475 ;
      RECT 90.8375 0.265 90.9025 0.415 ;
      RECT 90.835 0.27 90.905 0.41 ;
      RECT 89.8875 1.0425 89.9525 1.2825 ;
      RECT 89.885 1.095 89.955 1.235 ;
      RECT 89.7025 0.6575 89.7675 0.7925 ;
      RECT 89.045 0.6475 89.11 0.7825 ;
      RECT 89.045 0.685 89.7675 0.75 ;
      RECT 89.23 0.265 89.295 0.415 ;
      RECT 89.2275 0.27 89.2975 0.41 ;
      RECT 88.4 0.265 88.465 1.285 ;
      RECT 88.4 0.7875 88.695 0.8525 ;
      RECT 86.98 1.0425 87.045 1.2825 ;
      RECT 86.9775 1.095 87.0475 1.235 ;
      RECT 86.795 0.6575 86.86 0.7925 ;
      RECT 86.1375 0.6475 86.2025 0.7825 ;
      RECT 86.1375 0.685 86.86 0.75 ;
      RECT 86.3225 0.265 86.3875 0.415 ;
      RECT 86.32 0.27 86.39 0.41 ;
      RECT 85.4925 0.265 85.5575 1.285 ;
      RECT 85.4925 0.7875 85.7875 0.8525 ;
      RECT 84.0725 1.0425 84.1375 1.2825 ;
      RECT 84.07 1.095 84.14 1.235 ;
      RECT 83.8875 0.6575 83.9525 0.7925 ;
      RECT 83.23 0.6475 83.295 0.7825 ;
      RECT 83.23 0.685 83.9525 0.75 ;
      RECT 83.415 0.265 83.48 0.415 ;
      RECT 83.4125 0.27 83.4825 0.41 ;
      RECT 82.585 0.265 82.65 1.285 ;
      RECT 82.585 0.7875 82.88 0.8525 ;
      RECT 81.165 1.0425 81.23 1.2825 ;
      RECT 81.1625 1.095 81.2325 1.235 ;
      RECT 80.98 0.6575 81.045 0.7925 ;
      RECT 80.3225 0.6475 80.3875 0.7825 ;
      RECT 80.3225 0.685 81.045 0.75 ;
      RECT 80.5075 0.265 80.5725 0.415 ;
      RECT 80.505 0.27 80.575 0.41 ;
      RECT 79.6775 0.265 79.7425 1.285 ;
      RECT 79.6775 0.7875 79.9725 0.8525 ;
      RECT 78.2575 1.0425 78.3225 1.2825 ;
      RECT 78.255 1.095 78.325 1.235 ;
      RECT 78.0725 0.6575 78.1375 0.7925 ;
      RECT 77.415 0.6475 77.48 0.7825 ;
      RECT 77.415 0.685 78.1375 0.75 ;
      RECT 77.6 0.265 77.665 0.415 ;
      RECT 77.5975 0.27 77.6675 0.41 ;
      RECT 76.77 0.265 76.835 1.285 ;
      RECT 76.77 0.7875 77.065 0.8525 ;
      RECT 75.35 1.0425 75.415 1.2825 ;
      RECT 75.3475 1.095 75.4175 1.235 ;
      RECT 75.165 0.6575 75.23 0.7925 ;
      RECT 74.5075 0.6475 74.5725 0.7825 ;
      RECT 74.5075 0.685 75.23 0.75 ;
      RECT 74.6925 0.265 74.7575 0.415 ;
      RECT 74.69 0.27 74.76 0.41 ;
      RECT 73.8625 0.265 73.9275 1.285 ;
      RECT 73.8625 0.7875 74.1575 0.8525 ;
      RECT 72.4425 1.0425 72.5075 1.2825 ;
      RECT 72.44 1.095 72.51 1.235 ;
      RECT 72.2575 0.6575 72.3225 0.7925 ;
      RECT 71.6 0.6475 71.665 0.7825 ;
      RECT 71.6 0.685 72.3225 0.75 ;
      RECT 71.785 0.265 71.85 0.415 ;
      RECT 71.7825 0.27 71.8525 0.41 ;
      RECT 70.955 0.265 71.02 1.285 ;
      RECT 70.955 0.7875 71.25 0.8525 ;
      RECT 69.535 1.0425 69.6 1.2825 ;
      RECT 69.5325 1.095 69.6025 1.235 ;
      RECT 69.35 0.6575 69.415 0.7925 ;
      RECT 68.6925 0.6475 68.7575 0.7825 ;
      RECT 68.6925 0.685 69.415 0.75 ;
      RECT 68.8775 0.265 68.9425 0.415 ;
      RECT 68.875 0.27 68.945 0.41 ;
      RECT 68.0475 0.265 68.1125 1.285 ;
      RECT 68.0475 0.7875 68.3425 0.8525 ;
      RECT 66.6275 1.0425 66.6925 1.2825 ;
      RECT 66.625 1.095 66.695 1.235 ;
      RECT 66.4425 0.6575 66.5075 0.7925 ;
      RECT 65.785 0.6475 65.85 0.7825 ;
      RECT 65.785 0.685 66.5075 0.75 ;
      RECT 65.97 0.265 66.035 0.415 ;
      RECT 65.9675 0.27 66.0375 0.41 ;
      RECT 65.14 0.265 65.205 1.285 ;
      RECT 65.14 0.7875 65.435 0.8525 ;
      RECT 63.72 1.0425 63.785 1.2825 ;
      RECT 63.7175 1.095 63.7875 1.235 ;
      RECT 63.535 0.6575 63.6 0.7925 ;
      RECT 62.8775 0.6475 62.9425 0.7825 ;
      RECT 62.8775 0.685 63.6 0.75 ;
      RECT 63.0625 0.265 63.1275 0.415 ;
      RECT 63.06 0.27 63.13 0.41 ;
      RECT 62.2325 0.265 62.2975 1.285 ;
      RECT 62.2325 0.7875 62.5275 0.8525 ;
      RECT 60.8125 1.0425 60.8775 1.2825 ;
      RECT 60.81 1.095 60.88 1.235 ;
      RECT 60.6275 0.6575 60.6925 0.7925 ;
      RECT 59.97 0.6475 60.035 0.7825 ;
      RECT 59.97 0.685 60.6925 0.75 ;
      RECT 60.155 0.265 60.22 0.415 ;
      RECT 60.1525 0.27 60.2225 0.41 ;
      RECT 59.325 0.265 59.39 1.285 ;
      RECT 59.325 0.7875 59.62 0.8525 ;
      RECT 57.905 1.0425 57.97 1.2825 ;
      RECT 57.9025 1.095 57.9725 1.235 ;
      RECT 57.72 0.6575 57.785 0.7925 ;
      RECT 57.0625 0.6475 57.1275 0.7825 ;
      RECT 57.0625 0.685 57.785 0.75 ;
      RECT 57.2475 0.265 57.3125 0.415 ;
      RECT 57.245 0.27 57.315 0.41 ;
      RECT 56.4175 0.265 56.4825 1.285 ;
      RECT 56.4175 0.7875 56.7125 0.8525 ;
      RECT 54.9975 1.0425 55.0625 1.2825 ;
      RECT 54.995 1.095 55.065 1.235 ;
      RECT 54.8125 0.6575 54.8775 0.7925 ;
      RECT 54.155 0.6475 54.22 0.7825 ;
      RECT 54.155 0.685 54.8775 0.75 ;
      RECT 54.34 0.265 54.405 0.415 ;
      RECT 54.3375 0.27 54.4075 0.41 ;
      RECT 53.51 0.265 53.575 1.285 ;
      RECT 53.51 0.7875 53.805 0.8525 ;
      RECT 52.09 1.0425 52.155 1.2825 ;
      RECT 52.0875 1.095 52.1575 1.235 ;
      RECT 51.905 0.6575 51.97 0.7925 ;
      RECT 51.2475 0.6475 51.3125 0.7825 ;
      RECT 51.2475 0.685 51.97 0.75 ;
      RECT 51.4325 0.265 51.4975 0.415 ;
      RECT 51.43 0.27 51.5 0.41 ;
      RECT 50.6025 0.265 50.6675 1.285 ;
      RECT 50.6025 0.7875 50.8975 0.8525 ;
      RECT 49.1825 1.0425 49.2475 1.2825 ;
      RECT 49.18 1.095 49.25 1.235 ;
      RECT 48.9975 0.6575 49.0625 0.7925 ;
      RECT 48.34 0.6475 48.405 0.7825 ;
      RECT 48.34 0.685 49.0625 0.75 ;
      RECT 48.525 0.265 48.59 0.415 ;
      RECT 48.5225 0.27 48.5925 0.41 ;
      RECT 47.695 0.265 47.76 1.285 ;
      RECT 47.695 0.7875 47.99 0.8525 ;
      RECT 46.275 1.0425 46.34 1.2825 ;
      RECT 46.2725 1.095 46.3425 1.235 ;
      RECT 46.09 0.6575 46.155 0.7925 ;
      RECT 45.4325 0.6475 45.4975 0.7825 ;
      RECT 45.4325 0.685 46.155 0.75 ;
      RECT 45.6175 0.265 45.6825 0.415 ;
      RECT 45.615 0.27 45.685 0.41 ;
      RECT 44.7875 0.265 44.8525 1.285 ;
      RECT 44.7875 0.7875 45.0825 0.8525 ;
      RECT 43.3675 1.0425 43.4325 1.2825 ;
      RECT 43.365 1.095 43.435 1.235 ;
      RECT 43.1825 0.6575 43.2475 0.7925 ;
      RECT 42.525 0.6475 42.59 0.7825 ;
      RECT 42.525 0.685 43.2475 0.75 ;
      RECT 42.71 0.265 42.775 0.415 ;
      RECT 42.7075 0.27 42.7775 0.41 ;
      RECT 41.88 0.265 41.945 1.285 ;
      RECT 41.88 0.7875 42.175 0.8525 ;
      RECT 40.46 1.0425 40.525 1.2825 ;
      RECT 40.4575 1.095 40.5275 1.235 ;
      RECT 40.275 0.6575 40.34 0.7925 ;
      RECT 39.6175 0.6475 39.6825 0.7825 ;
      RECT 39.6175 0.685 40.34 0.75 ;
      RECT 39.8025 0.265 39.8675 0.415 ;
      RECT 39.8 0.27 39.87 0.41 ;
      RECT 38.9725 0.265 39.0375 1.285 ;
      RECT 38.9725 0.7875 39.2675 0.8525 ;
      RECT 37.5525 1.0425 37.6175 1.2825 ;
      RECT 37.55 1.095 37.62 1.235 ;
      RECT 37.3675 0.6575 37.4325 0.7925 ;
      RECT 36.71 0.6475 36.775 0.7825 ;
      RECT 36.71 0.685 37.4325 0.75 ;
      RECT 36.895 0.265 36.96 0.415 ;
      RECT 36.8925 0.27 36.9625 0.41 ;
      RECT 36.065 0.265 36.13 1.285 ;
      RECT 36.065 0.7875 36.36 0.8525 ;
      RECT 34.645 1.0425 34.71 1.2825 ;
      RECT 34.6425 1.095 34.7125 1.235 ;
      RECT 34.46 0.6575 34.525 0.7925 ;
      RECT 33.8025 0.6475 33.8675 0.7825 ;
      RECT 33.8025 0.685 34.525 0.75 ;
      RECT 33.9875 0.265 34.0525 0.415 ;
      RECT 33.985 0.27 34.055 0.41 ;
      RECT 33.1575 0.265 33.2225 1.285 ;
      RECT 33.1575 0.7875 33.4525 0.8525 ;
      RECT 31.7375 1.0425 31.8025 1.2825 ;
      RECT 31.735 1.095 31.805 1.235 ;
      RECT 31.5525 0.6575 31.6175 0.7925 ;
      RECT 30.895 0.6475 30.96 0.7825 ;
      RECT 30.895 0.685 31.6175 0.75 ;
      RECT 31.08 0.265 31.145 0.415 ;
      RECT 31.0775 0.27 31.1475 0.41 ;
      RECT 30.25 0.265 30.315 1.285 ;
      RECT 30.25 0.7875 30.545 0.8525 ;
      RECT 28.83 1.0425 28.895 1.2825 ;
      RECT 28.8275 1.095 28.8975 1.235 ;
      RECT 28.645 0.6575 28.71 0.7925 ;
      RECT 27.9875 0.6475 28.0525 0.7825 ;
      RECT 27.9875 0.685 28.71 0.75 ;
      RECT 28.1725 0.265 28.2375 0.415 ;
      RECT 28.17 0.27 28.24 0.41 ;
      RECT 27.3425 0.265 27.4075 1.285 ;
      RECT 27.3425 0.7875 27.6375 0.8525 ;
      RECT 25.9225 1.0425 25.9875 1.2825 ;
      RECT 25.92 1.095 25.99 1.235 ;
      RECT 25.7375 0.6575 25.8025 0.7925 ;
      RECT 25.08 0.6475 25.145 0.7825 ;
      RECT 25.08 0.685 25.8025 0.75 ;
      RECT 25.265 0.265 25.33 0.415 ;
      RECT 25.2625 0.27 25.3325 0.41 ;
      RECT 24.435 0.265 24.5 1.285 ;
      RECT 24.435 0.7875 24.73 0.8525 ;
      RECT 23.015 1.0425 23.08 1.2825 ;
      RECT 23.0125 1.095 23.0825 1.235 ;
      RECT 22.83 0.6575 22.895 0.7925 ;
      RECT 22.1725 0.6475 22.2375 0.7825 ;
      RECT 22.1725 0.685 22.895 0.75 ;
      RECT 22.3575 0.265 22.4225 0.415 ;
      RECT 22.355 0.27 22.425 0.41 ;
      RECT 21.5275 0.265 21.5925 1.285 ;
      RECT 21.5275 0.7875 21.8225 0.8525 ;
      RECT 20.1075 1.0425 20.1725 1.2825 ;
      RECT 20.105 1.095 20.175 1.235 ;
      RECT 19.9225 0.6575 19.9875 0.7925 ;
      RECT 19.265 0.6475 19.33 0.7825 ;
      RECT 19.265 0.685 19.9875 0.75 ;
      RECT 19.45 0.265 19.515 0.415 ;
      RECT 19.4475 0.27 19.5175 0.41 ;
      RECT 18.62 0.265 18.685 1.285 ;
      RECT 18.62 0.7875 18.915 0.8525 ;
      RECT 17.2 1.0425 17.265 1.2825 ;
      RECT 17.1975 1.095 17.2675 1.235 ;
      RECT 17.015 0.6575 17.08 0.7925 ;
      RECT 16.3575 0.6475 16.4225 0.7825 ;
      RECT 16.3575 0.685 17.08 0.75 ;
      RECT 16.5425 0.265 16.6075 0.415 ;
      RECT 16.54 0.27 16.61 0.41 ;
      RECT 15.7125 0.265 15.7775 1.285 ;
      RECT 15.7125 0.7875 16.0075 0.8525 ;
      RECT 14.2925 1.0425 14.3575 1.2825 ;
      RECT 14.29 1.095 14.36 1.235 ;
      RECT 14.1075 0.6575 14.1725 0.7925 ;
      RECT 13.45 0.6475 13.515 0.7825 ;
      RECT 13.45 0.685 14.1725 0.75 ;
      RECT 13.635 0.265 13.7 0.415 ;
      RECT 13.6325 0.27 13.7025 0.41 ;
      RECT 12.805 0.265 12.87 1.285 ;
      RECT 12.805 0.7875 13.1 0.8525 ;
      RECT 11.385 1.0425 11.45 1.2825 ;
      RECT 11.3825 1.095 11.4525 1.235 ;
      RECT 11.2 0.6575 11.265 0.7925 ;
      RECT 10.5425 0.6475 10.6075 0.7825 ;
      RECT 10.5425 0.685 11.265 0.75 ;
      RECT 10.7275 0.265 10.7925 0.415 ;
      RECT 10.725 0.27 10.795 0.41 ;
      RECT 9.8975 0.265 9.9625 1.285 ;
      RECT 9.8975 0.7875 10.1925 0.8525 ;
      RECT 8.4775 1.0425 8.5425 1.2825 ;
      RECT 8.475 1.095 8.545 1.235 ;
      RECT 8.2925 0.6575 8.3575 0.7925 ;
      RECT 7.635 0.6475 7.7 0.7825 ;
      RECT 7.635 0.685 8.3575 0.75 ;
      RECT 7.82 0.265 7.885 0.415 ;
      RECT 7.8175 0.27 7.8875 0.41 ;
      RECT 6.99 0.265 7.055 1.285 ;
      RECT 6.99 0.7875 7.285 0.8525 ;
      RECT 5.57 1.0425 5.635 1.2825 ;
      RECT 5.5675 1.095 5.6375 1.235 ;
      RECT 5.385 0.6575 5.45 0.7925 ;
      RECT 4.7275 0.6475 4.7925 0.7825 ;
      RECT 4.7275 0.685 5.45 0.75 ;
      RECT 4.9125 0.265 4.9775 0.415 ;
      RECT 4.91 0.27 4.98 0.41 ;
      RECT 4.0825 0.265 4.1475 1.285 ;
      RECT 4.0825 0.7875 4.3775 0.8525 ;
      RECT 2.6625 1.0425 2.7275 1.2825 ;
      RECT 2.66 1.095 2.73 1.235 ;
      RECT 2.4775 0.6575 2.5425 0.7925 ;
      RECT 1.82 0.6475 1.885 0.7825 ;
      RECT 1.82 0.685 2.5425 0.75 ;
      RECT 2.005 0.265 2.07 0.415 ;
      RECT 2.0025 0.27 2.0725 0.41 ;
      RECT 1.175 0.265 1.24 1.285 ;
      RECT 1.175 0.7875 1.47 0.8525 ;
      RECT 95.535 0.785 95.6 0.92 ;
      RECT 95.2975 0.2725 95.3625 0.4075 ;
      RECT 95.2975 1.0975 95.3625 1.2325 ;
      RECT 95.105 0.2725 95.17 0.4075 ;
      RECT 95.105 1.0975 95.17 1.2325 ;
      RECT 94.915 0.2725 94.98 0.4075 ;
      RECT 94.915 1.0975 94.98 1.2325 ;
      RECT 94.715 0.7075 94.78 0.8425 ;
      RECT 93.8575 0.75 93.9275 0.89 ;
      RECT 93.505 0.785 93.57 0.92 ;
      RECT 93.2675 0.2725 93.3325 0.4075 ;
      RECT 93.2675 1.0975 93.3325 1.2325 ;
      RECT 93.075 0.2725 93.14 0.4075 ;
      RECT 93.075 1.0975 93.14 1.2325 ;
      RECT 92.885 0.2725 92.95 0.4075 ;
      RECT 92.885 1.0975 92.95 1.2325 ;
      RECT 92.685 0.7075 92.75 0.8425 ;
      RECT 91.8275 0.75 91.8975 0.89 ;
      RECT 91.495 0.265 91.56 0.415 ;
      RECT 91.31 0.265 91.375 0.415 ;
      RECT 91.31 1.0425 91.375 1.2825 ;
      RECT 90.8375 1.0425 90.9025 1.2825 ;
      RECT 90.6525 0.265 90.7175 0.415 ;
      RECT 90.6525 1.0425 90.7175 1.2825 ;
      RECT 89.8875 0.265 89.9525 0.415 ;
      RECT 89.7025 0.265 89.7675 0.415 ;
      RECT 89.7025 1.0425 89.7675 1.2825 ;
      RECT 89.23 1.0425 89.295 1.2825 ;
      RECT 89.045 0.265 89.11 0.415 ;
      RECT 89.045 1.0425 89.11 1.2825 ;
      RECT 88.77 0.265 88.835 1.285 ;
      RECT 88.245 0.84 88.31 0.975 ;
      RECT 87.9375 0.265 88.0025 0.415 ;
      RECT 87.9375 1.0425 88.0025 1.2825 ;
      RECT 87.7525 0.265 87.8175 0.415 ;
      RECT 87.7525 1.0425 87.8175 1.2825 ;
      RECT 87.5675 0.265 87.6325 0.415 ;
      RECT 87.5675 1.0425 87.6325 1.2825 ;
      RECT 86.98 0.265 87.045 0.415 ;
      RECT 86.795 0.265 86.86 0.415 ;
      RECT 86.795 1.0425 86.86 1.2825 ;
      RECT 86.3225 1.0425 86.3875 1.2825 ;
      RECT 86.1375 0.265 86.2025 0.415 ;
      RECT 86.1375 1.0425 86.2025 1.2825 ;
      RECT 85.8625 0.265 85.9275 1.285 ;
      RECT 85.3375 0.84 85.4025 0.975 ;
      RECT 85.03 0.265 85.095 0.415 ;
      RECT 85.03 1.0425 85.095 1.2825 ;
      RECT 84.845 0.265 84.91 0.415 ;
      RECT 84.845 1.0425 84.91 1.2825 ;
      RECT 84.66 0.265 84.725 0.415 ;
      RECT 84.66 1.0425 84.725 1.2825 ;
      RECT 84.0725 0.265 84.1375 0.415 ;
      RECT 83.8875 0.265 83.9525 0.415 ;
      RECT 83.8875 1.0425 83.9525 1.2825 ;
      RECT 83.415 1.0425 83.48 1.2825 ;
      RECT 83.23 0.265 83.295 0.415 ;
      RECT 83.23 1.0425 83.295 1.2825 ;
      RECT 82.955 0.265 83.02 1.285 ;
      RECT 82.43 0.84 82.495 0.975 ;
      RECT 82.1225 0.265 82.1875 0.415 ;
      RECT 82.1225 1.0425 82.1875 1.2825 ;
      RECT 81.9375 0.265 82.0025 0.415 ;
      RECT 81.9375 1.0425 82.0025 1.2825 ;
      RECT 81.7525 0.265 81.8175 0.415 ;
      RECT 81.7525 1.0425 81.8175 1.2825 ;
      RECT 81.165 0.265 81.23 0.415 ;
      RECT 80.98 0.265 81.045 0.415 ;
      RECT 80.98 1.0425 81.045 1.2825 ;
      RECT 80.5075 1.0425 80.5725 1.2825 ;
      RECT 80.3225 0.265 80.3875 0.415 ;
      RECT 80.3225 1.0425 80.3875 1.2825 ;
      RECT 80.0475 0.265 80.1125 1.285 ;
      RECT 79.5225 0.84 79.5875 0.975 ;
      RECT 79.215 0.265 79.28 0.415 ;
      RECT 79.215 1.0425 79.28 1.2825 ;
      RECT 79.03 0.265 79.095 0.415 ;
      RECT 79.03 1.0425 79.095 1.2825 ;
      RECT 78.845 0.265 78.91 0.415 ;
      RECT 78.845 1.0425 78.91 1.2825 ;
      RECT 78.2575 0.265 78.3225 0.415 ;
      RECT 78.0725 0.265 78.1375 0.415 ;
      RECT 78.0725 1.0425 78.1375 1.2825 ;
      RECT 77.6 1.0425 77.665 1.2825 ;
      RECT 77.415 0.265 77.48 0.415 ;
      RECT 77.415 1.0425 77.48 1.2825 ;
      RECT 77.14 0.265 77.205 1.285 ;
      RECT 76.615 0.84 76.68 0.975 ;
      RECT 76.3075 0.265 76.3725 0.415 ;
      RECT 76.3075 1.0425 76.3725 1.2825 ;
      RECT 76.1225 0.265 76.1875 0.415 ;
      RECT 76.1225 1.0425 76.1875 1.2825 ;
      RECT 75.9375 0.265 76.0025 0.415 ;
      RECT 75.9375 1.0425 76.0025 1.2825 ;
      RECT 75.35 0.265 75.415 0.415 ;
      RECT 75.165 0.265 75.23 0.415 ;
      RECT 75.165 1.0425 75.23 1.2825 ;
      RECT 74.6925 1.0425 74.7575 1.2825 ;
      RECT 74.5075 0.265 74.5725 0.415 ;
      RECT 74.5075 1.0425 74.5725 1.2825 ;
      RECT 74.2325 0.265 74.2975 1.285 ;
      RECT 73.7075 0.84 73.7725 0.975 ;
      RECT 73.4 0.265 73.465 0.415 ;
      RECT 73.4 1.0425 73.465 1.2825 ;
      RECT 73.215 0.265 73.28 0.415 ;
      RECT 73.215 1.0425 73.28 1.2825 ;
      RECT 73.03 0.265 73.095 0.415 ;
      RECT 73.03 1.0425 73.095 1.2825 ;
      RECT 72.4425 0.265 72.5075 0.415 ;
      RECT 72.2575 0.265 72.3225 0.415 ;
      RECT 72.2575 1.0425 72.3225 1.2825 ;
      RECT 71.785 1.0425 71.85 1.2825 ;
      RECT 71.6 0.265 71.665 0.415 ;
      RECT 71.6 1.0425 71.665 1.2825 ;
      RECT 71.325 0.265 71.39 1.285 ;
      RECT 70.8 0.84 70.865 0.975 ;
      RECT 70.4925 0.265 70.5575 0.415 ;
      RECT 70.4925 1.0425 70.5575 1.2825 ;
      RECT 70.3075 0.265 70.3725 0.415 ;
      RECT 70.3075 1.0425 70.3725 1.2825 ;
      RECT 70.1225 0.265 70.1875 0.415 ;
      RECT 70.1225 1.0425 70.1875 1.2825 ;
      RECT 69.535 0.265 69.6 0.415 ;
      RECT 69.35 0.265 69.415 0.415 ;
      RECT 69.35 1.0425 69.415 1.2825 ;
      RECT 68.8775 1.0425 68.9425 1.2825 ;
      RECT 68.6925 0.265 68.7575 0.415 ;
      RECT 68.6925 1.0425 68.7575 1.2825 ;
      RECT 68.4175 0.265 68.4825 1.285 ;
      RECT 67.8925 0.84 67.9575 0.975 ;
      RECT 67.585 0.265 67.65 0.415 ;
      RECT 67.585 1.0425 67.65 1.2825 ;
      RECT 67.4 0.265 67.465 0.415 ;
      RECT 67.4 1.0425 67.465 1.2825 ;
      RECT 67.215 0.265 67.28 0.415 ;
      RECT 67.215 1.0425 67.28 1.2825 ;
      RECT 66.6275 0.265 66.6925 0.415 ;
      RECT 66.4425 0.265 66.5075 0.415 ;
      RECT 66.4425 1.0425 66.5075 1.2825 ;
      RECT 65.97 1.0425 66.035 1.2825 ;
      RECT 65.785 0.265 65.85 0.415 ;
      RECT 65.785 1.0425 65.85 1.2825 ;
      RECT 65.51 0.265 65.575 1.285 ;
      RECT 64.985 0.84 65.05 0.975 ;
      RECT 64.6775 0.265 64.7425 0.415 ;
      RECT 64.6775 1.0425 64.7425 1.2825 ;
      RECT 64.4925 0.265 64.5575 0.415 ;
      RECT 64.4925 1.0425 64.5575 1.2825 ;
      RECT 64.3075 0.265 64.3725 0.415 ;
      RECT 64.3075 1.0425 64.3725 1.2825 ;
      RECT 63.72 0.265 63.785 0.415 ;
      RECT 63.535 0.265 63.6 0.415 ;
      RECT 63.535 1.0425 63.6 1.2825 ;
      RECT 63.0625 1.0425 63.1275 1.2825 ;
      RECT 62.8775 0.265 62.9425 0.415 ;
      RECT 62.8775 1.0425 62.9425 1.2825 ;
      RECT 62.6025 0.265 62.6675 1.285 ;
      RECT 62.0775 0.84 62.1425 0.975 ;
      RECT 61.77 0.265 61.835 0.415 ;
      RECT 61.77 1.0425 61.835 1.2825 ;
      RECT 61.585 0.265 61.65 0.415 ;
      RECT 61.585 1.0425 61.65 1.2825 ;
      RECT 61.4 0.265 61.465 0.415 ;
      RECT 61.4 1.0425 61.465 1.2825 ;
      RECT 60.8125 0.265 60.8775 0.415 ;
      RECT 60.6275 0.265 60.6925 0.415 ;
      RECT 60.6275 1.0425 60.6925 1.2825 ;
      RECT 60.155 1.0425 60.22 1.2825 ;
      RECT 59.97 0.265 60.035 0.415 ;
      RECT 59.97 1.0425 60.035 1.2825 ;
      RECT 59.695 0.265 59.76 1.285 ;
      RECT 59.17 0.84 59.235 0.975 ;
      RECT 58.8625 0.265 58.9275 0.415 ;
      RECT 58.8625 1.0425 58.9275 1.2825 ;
      RECT 58.6775 0.265 58.7425 0.415 ;
      RECT 58.6775 1.0425 58.7425 1.2825 ;
      RECT 58.4925 0.265 58.5575 0.415 ;
      RECT 58.4925 1.0425 58.5575 1.2825 ;
      RECT 57.905 0.265 57.97 0.415 ;
      RECT 57.72 0.265 57.785 0.415 ;
      RECT 57.72 1.0425 57.785 1.2825 ;
      RECT 57.2475 1.0425 57.3125 1.2825 ;
      RECT 57.0625 0.265 57.1275 0.415 ;
      RECT 57.0625 1.0425 57.1275 1.2825 ;
      RECT 56.7875 0.265 56.8525 1.285 ;
      RECT 56.2625 0.84 56.3275 0.975 ;
      RECT 55.955 0.265 56.02 0.415 ;
      RECT 55.955 1.0425 56.02 1.2825 ;
      RECT 55.77 0.265 55.835 0.415 ;
      RECT 55.77 1.0425 55.835 1.2825 ;
      RECT 55.585 0.265 55.65 0.415 ;
      RECT 55.585 1.0425 55.65 1.2825 ;
      RECT 54.9975 0.265 55.0625 0.415 ;
      RECT 54.8125 0.265 54.8775 0.415 ;
      RECT 54.8125 1.0425 54.8775 1.2825 ;
      RECT 54.34 1.0425 54.405 1.2825 ;
      RECT 54.155 0.265 54.22 0.415 ;
      RECT 54.155 1.0425 54.22 1.2825 ;
      RECT 53.88 0.265 53.945 1.285 ;
      RECT 53.355 0.84 53.42 0.975 ;
      RECT 53.0475 0.265 53.1125 0.415 ;
      RECT 53.0475 1.0425 53.1125 1.2825 ;
      RECT 52.8625 0.265 52.9275 0.415 ;
      RECT 52.8625 1.0425 52.9275 1.2825 ;
      RECT 52.6775 0.265 52.7425 0.415 ;
      RECT 52.6775 1.0425 52.7425 1.2825 ;
      RECT 52.09 0.265 52.155 0.415 ;
      RECT 51.905 0.265 51.97 0.415 ;
      RECT 51.905 1.0425 51.97 1.2825 ;
      RECT 51.4325 1.0425 51.4975 1.2825 ;
      RECT 51.2475 0.265 51.3125 0.415 ;
      RECT 51.2475 1.0425 51.3125 1.2825 ;
      RECT 50.9725 0.265 51.0375 1.285 ;
      RECT 50.4475 0.84 50.5125 0.975 ;
      RECT 50.14 0.265 50.205 0.415 ;
      RECT 50.14 1.0425 50.205 1.2825 ;
      RECT 49.955 0.265 50.02 0.415 ;
      RECT 49.955 1.0425 50.02 1.2825 ;
      RECT 49.77 0.265 49.835 0.415 ;
      RECT 49.77 1.0425 49.835 1.2825 ;
      RECT 49.1825 0.265 49.2475 0.415 ;
      RECT 48.9975 0.265 49.0625 0.415 ;
      RECT 48.9975 1.0425 49.0625 1.2825 ;
      RECT 48.525 1.0425 48.59 1.2825 ;
      RECT 48.34 0.265 48.405 0.415 ;
      RECT 48.34 1.0425 48.405 1.2825 ;
      RECT 48.065 0.265 48.13 1.285 ;
      RECT 47.54 0.84 47.605 0.975 ;
      RECT 47.2325 0.265 47.2975 0.415 ;
      RECT 47.2325 1.0425 47.2975 1.2825 ;
      RECT 47.0475 0.265 47.1125 0.415 ;
      RECT 47.0475 1.0425 47.1125 1.2825 ;
      RECT 46.8625 0.265 46.9275 0.415 ;
      RECT 46.8625 1.0425 46.9275 1.2825 ;
      RECT 46.275 0.265 46.34 0.415 ;
      RECT 46.09 0.265 46.155 0.415 ;
      RECT 46.09 1.0425 46.155 1.2825 ;
      RECT 45.6175 1.0425 45.6825 1.2825 ;
      RECT 45.4325 0.265 45.4975 0.415 ;
      RECT 45.4325 1.0425 45.4975 1.2825 ;
      RECT 45.1575 0.265 45.2225 1.285 ;
      RECT 44.6325 0.84 44.6975 0.975 ;
      RECT 44.325 0.265 44.39 0.415 ;
      RECT 44.325 1.0425 44.39 1.2825 ;
      RECT 44.14 0.265 44.205 0.415 ;
      RECT 44.14 1.0425 44.205 1.2825 ;
      RECT 43.955 0.265 44.02 0.415 ;
      RECT 43.955 1.0425 44.02 1.2825 ;
      RECT 43.3675 0.265 43.4325 0.415 ;
      RECT 43.1825 0.265 43.2475 0.415 ;
      RECT 43.1825 1.0425 43.2475 1.2825 ;
      RECT 42.71 1.0425 42.775 1.2825 ;
      RECT 42.525 0.265 42.59 0.415 ;
      RECT 42.525 1.0425 42.59 1.2825 ;
      RECT 42.25 0.265 42.315 1.285 ;
      RECT 41.725 0.84 41.79 0.975 ;
      RECT 41.4175 0.265 41.4825 0.415 ;
      RECT 41.4175 1.0425 41.4825 1.2825 ;
      RECT 41.2325 0.265 41.2975 0.415 ;
      RECT 41.2325 1.0425 41.2975 1.2825 ;
      RECT 41.0475 0.265 41.1125 0.415 ;
      RECT 41.0475 1.0425 41.1125 1.2825 ;
      RECT 40.46 0.265 40.525 0.415 ;
      RECT 40.275 0.265 40.34 0.415 ;
      RECT 40.275 1.0425 40.34 1.2825 ;
      RECT 39.8025 1.0425 39.8675 1.2825 ;
      RECT 39.6175 0.265 39.6825 0.415 ;
      RECT 39.6175 1.0425 39.6825 1.2825 ;
      RECT 39.3425 0.265 39.4075 1.285 ;
      RECT 38.8175 0.84 38.8825 0.975 ;
      RECT 38.51 0.265 38.575 0.415 ;
      RECT 38.51 1.0425 38.575 1.2825 ;
      RECT 38.325 0.265 38.39 0.415 ;
      RECT 38.325 1.0425 38.39 1.2825 ;
      RECT 38.14 0.265 38.205 0.415 ;
      RECT 38.14 1.0425 38.205 1.2825 ;
      RECT 37.5525 0.265 37.6175 0.415 ;
      RECT 37.3675 0.265 37.4325 0.415 ;
      RECT 37.3675 1.0425 37.4325 1.2825 ;
      RECT 36.895 1.0425 36.96 1.2825 ;
      RECT 36.71 0.265 36.775 0.415 ;
      RECT 36.71 1.0425 36.775 1.2825 ;
      RECT 36.435 0.265 36.5 1.285 ;
      RECT 35.91 0.84 35.975 0.975 ;
      RECT 35.6025 0.265 35.6675 0.415 ;
      RECT 35.6025 1.0425 35.6675 1.2825 ;
      RECT 35.4175 0.265 35.4825 0.415 ;
      RECT 35.4175 1.0425 35.4825 1.2825 ;
      RECT 35.2325 0.265 35.2975 0.415 ;
      RECT 35.2325 1.0425 35.2975 1.2825 ;
      RECT 34.645 0.265 34.71 0.415 ;
      RECT 34.46 0.265 34.525 0.415 ;
      RECT 34.46 1.0425 34.525 1.2825 ;
      RECT 33.9875 1.0425 34.0525 1.2825 ;
      RECT 33.8025 0.265 33.8675 0.415 ;
      RECT 33.8025 1.0425 33.8675 1.2825 ;
      RECT 33.5275 0.265 33.5925 1.285 ;
      RECT 33.0025 0.84 33.0675 0.975 ;
      RECT 32.695 0.265 32.76 0.415 ;
      RECT 32.695 1.0425 32.76 1.2825 ;
      RECT 32.51 0.265 32.575 0.415 ;
      RECT 32.51 1.0425 32.575 1.2825 ;
      RECT 32.325 0.265 32.39 0.415 ;
      RECT 32.325 1.0425 32.39 1.2825 ;
      RECT 31.7375 0.265 31.8025 0.415 ;
      RECT 31.5525 0.265 31.6175 0.415 ;
      RECT 31.5525 1.0425 31.6175 1.2825 ;
      RECT 31.08 1.0425 31.145 1.2825 ;
      RECT 30.895 0.265 30.96 0.415 ;
      RECT 30.895 1.0425 30.96 1.2825 ;
      RECT 30.62 0.265 30.685 1.285 ;
      RECT 30.095 0.84 30.16 0.975 ;
      RECT 29.7875 0.265 29.8525 0.415 ;
      RECT 29.7875 1.0425 29.8525 1.2825 ;
      RECT 29.6025 0.265 29.6675 0.415 ;
      RECT 29.6025 1.0425 29.6675 1.2825 ;
      RECT 29.4175 0.265 29.4825 0.415 ;
      RECT 29.4175 1.0425 29.4825 1.2825 ;
      RECT 28.83 0.265 28.895 0.415 ;
      RECT 28.645 0.265 28.71 0.415 ;
      RECT 28.645 1.0425 28.71 1.2825 ;
      RECT 28.1725 1.0425 28.2375 1.2825 ;
      RECT 27.9875 0.265 28.0525 0.415 ;
      RECT 27.9875 1.0425 28.0525 1.2825 ;
      RECT 27.7125 0.265 27.7775 1.285 ;
      RECT 27.1875 0.84 27.2525 0.975 ;
      RECT 26.88 0.265 26.945 0.415 ;
      RECT 26.88 1.0425 26.945 1.2825 ;
      RECT 26.695 0.265 26.76 0.415 ;
      RECT 26.695 1.0425 26.76 1.2825 ;
      RECT 26.51 0.265 26.575 0.415 ;
      RECT 26.51 1.0425 26.575 1.2825 ;
      RECT 25.9225 0.265 25.9875 0.415 ;
      RECT 25.7375 0.265 25.8025 0.415 ;
      RECT 25.7375 1.0425 25.8025 1.2825 ;
      RECT 25.265 1.0425 25.33 1.2825 ;
      RECT 25.08 0.265 25.145 0.415 ;
      RECT 25.08 1.0425 25.145 1.2825 ;
      RECT 24.805 0.265 24.87 1.285 ;
      RECT 24.28 0.84 24.345 0.975 ;
      RECT 23.9725 0.265 24.0375 0.415 ;
      RECT 23.9725 1.0425 24.0375 1.2825 ;
      RECT 23.7875 0.265 23.8525 0.415 ;
      RECT 23.7875 1.0425 23.8525 1.2825 ;
      RECT 23.6025 0.265 23.6675 0.415 ;
      RECT 23.6025 1.0425 23.6675 1.2825 ;
      RECT 23.015 0.265 23.08 0.415 ;
      RECT 22.83 0.265 22.895 0.415 ;
      RECT 22.83 1.0425 22.895 1.2825 ;
      RECT 22.3575 1.0425 22.4225 1.2825 ;
      RECT 22.1725 0.265 22.2375 0.415 ;
      RECT 22.1725 1.0425 22.2375 1.2825 ;
      RECT 21.8975 0.265 21.9625 1.285 ;
      RECT 21.3725 0.84 21.4375 0.975 ;
      RECT 21.065 0.265 21.13 0.415 ;
      RECT 21.065 1.0425 21.13 1.2825 ;
      RECT 20.88 0.265 20.945 0.415 ;
      RECT 20.88 1.0425 20.945 1.2825 ;
      RECT 20.695 0.265 20.76 0.415 ;
      RECT 20.695 1.0425 20.76 1.2825 ;
      RECT 20.1075 0.265 20.1725 0.415 ;
      RECT 19.9225 0.265 19.9875 0.415 ;
      RECT 19.9225 1.0425 19.9875 1.2825 ;
      RECT 19.45 1.0425 19.515 1.2825 ;
      RECT 19.265 0.265 19.33 0.415 ;
      RECT 19.265 1.0425 19.33 1.2825 ;
      RECT 18.99 0.265 19.055 1.285 ;
      RECT 18.465 0.84 18.53 0.975 ;
      RECT 18.1575 0.265 18.2225 0.415 ;
      RECT 18.1575 1.0425 18.2225 1.2825 ;
      RECT 17.9725 0.265 18.0375 0.415 ;
      RECT 17.9725 1.0425 18.0375 1.2825 ;
      RECT 17.7875 0.265 17.8525 0.415 ;
      RECT 17.7875 1.0425 17.8525 1.2825 ;
      RECT 17.2 0.265 17.265 0.415 ;
      RECT 17.015 0.265 17.08 0.415 ;
      RECT 17.015 1.0425 17.08 1.2825 ;
      RECT 16.5425 1.0425 16.6075 1.2825 ;
      RECT 16.3575 0.265 16.4225 0.415 ;
      RECT 16.3575 1.0425 16.4225 1.2825 ;
      RECT 16.0825 0.265 16.1475 1.285 ;
      RECT 15.5575 0.84 15.6225 0.975 ;
      RECT 15.25 0.265 15.315 0.415 ;
      RECT 15.25 1.0425 15.315 1.2825 ;
      RECT 15.065 0.265 15.13 0.415 ;
      RECT 15.065 1.0425 15.13 1.2825 ;
      RECT 14.88 0.265 14.945 0.415 ;
      RECT 14.88 1.0425 14.945 1.2825 ;
      RECT 14.2925 0.265 14.3575 0.415 ;
      RECT 14.1075 0.265 14.1725 0.415 ;
      RECT 14.1075 1.0425 14.1725 1.2825 ;
      RECT 13.635 1.0425 13.7 1.2825 ;
      RECT 13.45 0.265 13.515 0.415 ;
      RECT 13.45 1.0425 13.515 1.2825 ;
      RECT 13.175 0.265 13.24 1.285 ;
      RECT 12.65 0.84 12.715 0.975 ;
      RECT 12.3425 0.265 12.4075 0.415 ;
      RECT 12.3425 1.0425 12.4075 1.2825 ;
      RECT 12.1575 0.265 12.2225 0.415 ;
      RECT 12.1575 1.0425 12.2225 1.2825 ;
      RECT 11.9725 0.265 12.0375 0.415 ;
      RECT 11.9725 1.0425 12.0375 1.2825 ;
      RECT 11.385 0.265 11.45 0.415 ;
      RECT 11.2 0.265 11.265 0.415 ;
      RECT 11.2 1.0425 11.265 1.2825 ;
      RECT 10.7275 1.0425 10.7925 1.2825 ;
      RECT 10.5425 0.265 10.6075 0.415 ;
      RECT 10.5425 1.0425 10.6075 1.2825 ;
      RECT 10.2675 0.265 10.3325 1.285 ;
      RECT 9.7425 0.84 9.8075 0.975 ;
      RECT 9.435 0.265 9.5 0.415 ;
      RECT 9.435 1.0425 9.5 1.2825 ;
      RECT 9.25 0.265 9.315 0.415 ;
      RECT 9.25 1.0425 9.315 1.2825 ;
      RECT 9.065 0.265 9.13 0.415 ;
      RECT 9.065 1.0425 9.13 1.2825 ;
      RECT 8.4775 0.265 8.5425 0.415 ;
      RECT 8.2925 0.265 8.3575 0.415 ;
      RECT 8.2925 1.0425 8.3575 1.2825 ;
      RECT 7.82 1.0425 7.885 1.2825 ;
      RECT 7.635 0.265 7.7 0.415 ;
      RECT 7.635 1.0425 7.7 1.2825 ;
      RECT 7.36 0.265 7.425 1.285 ;
      RECT 6.835 0.84 6.9 0.975 ;
      RECT 6.5275 0.265 6.5925 0.415 ;
      RECT 6.5275 1.0425 6.5925 1.2825 ;
      RECT 6.3425 0.265 6.4075 0.415 ;
      RECT 6.3425 1.0425 6.4075 1.2825 ;
      RECT 6.1575 0.265 6.2225 0.415 ;
      RECT 6.1575 1.0425 6.2225 1.2825 ;
      RECT 5.57 0.265 5.635 0.415 ;
      RECT 5.385 0.265 5.45 0.415 ;
      RECT 5.385 1.0425 5.45 1.2825 ;
      RECT 4.9125 1.0425 4.9775 1.2825 ;
      RECT 4.7275 0.265 4.7925 0.415 ;
      RECT 4.7275 1.0425 4.7925 1.2825 ;
      RECT 4.4525 0.265 4.5175 1.285 ;
      RECT 3.9275 0.84 3.9925 0.975 ;
      RECT 3.62 0.265 3.685 0.415 ;
      RECT 3.62 1.0425 3.685 1.2825 ;
      RECT 3.435 0.265 3.5 0.415 ;
      RECT 3.435 1.0425 3.5 1.2825 ;
      RECT 3.25 0.265 3.315 0.415 ;
      RECT 3.25 1.0425 3.315 1.2825 ;
      RECT 2.6625 0.265 2.7275 0.415 ;
      RECT 2.4775 0.265 2.5425 0.415 ;
      RECT 2.4775 1.0425 2.5425 1.2825 ;
      RECT 2.005 1.0425 2.07 1.2825 ;
      RECT 1.82 0.265 1.885 0.415 ;
      RECT 1.82 1.0425 1.885 1.2825 ;
      RECT 1.545 0.265 1.61 1.285 ;
      RECT 1.02 0.84 1.085 0.975 ;
      RECT 0.7125 0.265 0.7775 0.415 ;
      RECT 0.7125 1.0425 0.7775 1.2825 ;
      RECT 0.5275 0.265 0.5925 0.415 ;
      RECT 0.5275 1.0425 0.5925 1.2825 ;
      RECT 0.3425 0.265 0.4075 0.415 ;
      RECT 0.3425 1.0425 0.4075 1.2825 ;
    LAYER metal2 ;
      RECT 95.1025 1.3075 95.6025 1.3775 ;
      RECT 95.5325 0.785 95.6025 1.3775 ;
      RECT 95.1025 0.265 95.1725 1.3775 ;
      RECT 94.7125 0.525 94.7825 0.8425 ;
      RECT 94.015 0.49 94.085 0.625 ;
      RECT 94.015 0.525 94.7825 0.595 ;
      RECT 93.0725 1.3075 93.5725 1.3775 ;
      RECT 93.5025 0.785 93.5725 1.3775 ;
      RECT 93.0725 0.265 93.1425 1.3775 ;
      RECT 92.6825 0.525 92.7525 0.8425 ;
      RECT 91.985 0.49 92.055 0.625 ;
      RECT 91.985 0.525 92.7525 0.595 ;
      RECT 89.0425 0.2725 89.1125 1.2325 ;
      RECT 88.3975 0.2725 88.4675 0.4075 ;
      RECT 88.3975 0.3075 89.1125 0.3775 ;
      RECT 87.935 0.2725 88.005 1.2325 ;
      RECT 88.7675 0.6225 88.8375 0.7575 ;
      RECT 87.935 0.665 88.8375 0.735 ;
      RECT 87.75 1.315 88.3125 1.385 ;
      RECT 88.2425 0.84 88.3125 1.385 ;
      RECT 87.75 0.2725 87.82 1.385 ;
      RECT 87.565 1.0975 87.635 1.2325 ;
      RECT 87.565 1.1325 87.82 1.2025 ;
      RECT 87.565 0.2725 87.635 0.4075 ;
      RECT 87.565 0.3075 87.82 0.3775 ;
      RECT 86.135 0.2725 86.205 1.2325 ;
      RECT 85.49 0.2725 85.56 0.4075 ;
      RECT 85.49 0.3075 86.205 0.3775 ;
      RECT 85.0275 0.2725 85.0975 1.2325 ;
      RECT 85.86 0.6225 85.93 0.7575 ;
      RECT 85.0275 0.665 85.93 0.735 ;
      RECT 84.8425 1.315 85.405 1.385 ;
      RECT 85.335 0.84 85.405 1.385 ;
      RECT 84.8425 0.2725 84.9125 1.385 ;
      RECT 84.6575 1.0975 84.7275 1.2325 ;
      RECT 84.6575 1.1325 84.9125 1.2025 ;
      RECT 84.6575 0.2725 84.7275 0.4075 ;
      RECT 84.6575 0.3075 84.9125 0.3775 ;
      RECT 83.2275 0.2725 83.2975 1.2325 ;
      RECT 82.5825 0.2725 82.6525 0.4075 ;
      RECT 82.5825 0.3075 83.2975 0.3775 ;
      RECT 82.12 0.2725 82.19 1.2325 ;
      RECT 82.9525 0.6225 83.0225 0.7575 ;
      RECT 82.12 0.665 83.0225 0.735 ;
      RECT 81.935 1.315 82.4975 1.385 ;
      RECT 82.4275 0.84 82.4975 1.385 ;
      RECT 81.935 0.2725 82.005 1.385 ;
      RECT 81.75 1.0975 81.82 1.2325 ;
      RECT 81.75 1.1325 82.005 1.2025 ;
      RECT 81.75 0.2725 81.82 0.4075 ;
      RECT 81.75 0.3075 82.005 0.3775 ;
      RECT 80.32 0.2725 80.39 1.2325 ;
      RECT 79.675 0.2725 79.745 0.4075 ;
      RECT 79.675 0.3075 80.39 0.3775 ;
      RECT 79.2125 0.2725 79.2825 1.2325 ;
      RECT 80.045 0.6225 80.115 0.7575 ;
      RECT 79.2125 0.665 80.115 0.735 ;
      RECT 79.0275 1.315 79.59 1.385 ;
      RECT 79.52 0.84 79.59 1.385 ;
      RECT 79.0275 0.2725 79.0975 1.385 ;
      RECT 78.8425 1.0975 78.9125 1.2325 ;
      RECT 78.8425 1.1325 79.0975 1.2025 ;
      RECT 78.8425 0.2725 78.9125 0.4075 ;
      RECT 78.8425 0.3075 79.0975 0.3775 ;
      RECT 77.4125 0.2725 77.4825 1.2325 ;
      RECT 76.7675 0.2725 76.8375 0.4075 ;
      RECT 76.7675 0.3075 77.4825 0.3775 ;
      RECT 76.305 0.2725 76.375 1.2325 ;
      RECT 77.1375 0.6225 77.2075 0.7575 ;
      RECT 76.305 0.665 77.2075 0.735 ;
      RECT 76.12 1.315 76.6825 1.385 ;
      RECT 76.6125 0.84 76.6825 1.385 ;
      RECT 76.12 0.2725 76.19 1.385 ;
      RECT 75.935 1.0975 76.005 1.2325 ;
      RECT 75.935 1.1325 76.19 1.2025 ;
      RECT 75.935 0.2725 76.005 0.4075 ;
      RECT 75.935 0.3075 76.19 0.3775 ;
      RECT 74.505 0.2725 74.575 1.2325 ;
      RECT 73.86 0.2725 73.93 0.4075 ;
      RECT 73.86 0.3075 74.575 0.3775 ;
      RECT 73.3975 0.2725 73.4675 1.2325 ;
      RECT 74.23 0.6225 74.3 0.7575 ;
      RECT 73.3975 0.665 74.3 0.735 ;
      RECT 73.2125 1.315 73.775 1.385 ;
      RECT 73.705 0.84 73.775 1.385 ;
      RECT 73.2125 0.2725 73.2825 1.385 ;
      RECT 73.0275 1.0975 73.0975 1.2325 ;
      RECT 73.0275 1.1325 73.2825 1.2025 ;
      RECT 73.0275 0.2725 73.0975 0.4075 ;
      RECT 73.0275 0.3075 73.2825 0.3775 ;
      RECT 71.5975 0.2725 71.6675 1.2325 ;
      RECT 70.9525 0.2725 71.0225 0.4075 ;
      RECT 70.9525 0.3075 71.6675 0.3775 ;
      RECT 70.49 0.2725 70.56 1.2325 ;
      RECT 71.3225 0.6225 71.3925 0.7575 ;
      RECT 70.49 0.665 71.3925 0.735 ;
      RECT 70.305 1.315 70.8675 1.385 ;
      RECT 70.7975 0.84 70.8675 1.385 ;
      RECT 70.305 0.2725 70.375 1.385 ;
      RECT 70.12 1.0975 70.19 1.2325 ;
      RECT 70.12 1.1325 70.375 1.2025 ;
      RECT 70.12 0.2725 70.19 0.4075 ;
      RECT 70.12 0.3075 70.375 0.3775 ;
      RECT 68.69 0.2725 68.76 1.2325 ;
      RECT 68.045 0.2725 68.115 0.4075 ;
      RECT 68.045 0.3075 68.76 0.3775 ;
      RECT 67.5825 0.2725 67.6525 1.2325 ;
      RECT 68.415 0.6225 68.485 0.7575 ;
      RECT 67.5825 0.665 68.485 0.735 ;
      RECT 67.3975 1.315 67.96 1.385 ;
      RECT 67.89 0.84 67.96 1.385 ;
      RECT 67.3975 0.2725 67.4675 1.385 ;
      RECT 67.2125 1.0975 67.2825 1.2325 ;
      RECT 67.2125 1.1325 67.4675 1.2025 ;
      RECT 67.2125 0.2725 67.2825 0.4075 ;
      RECT 67.2125 0.3075 67.4675 0.3775 ;
      RECT 65.7825 0.2725 65.8525 1.2325 ;
      RECT 65.1375 0.2725 65.2075 0.4075 ;
      RECT 65.1375 0.3075 65.8525 0.3775 ;
      RECT 64.675 0.2725 64.745 1.2325 ;
      RECT 65.5075 0.6225 65.5775 0.7575 ;
      RECT 64.675 0.665 65.5775 0.735 ;
      RECT 64.49 1.315 65.0525 1.385 ;
      RECT 64.9825 0.84 65.0525 1.385 ;
      RECT 64.49 0.2725 64.56 1.385 ;
      RECT 64.305 1.0975 64.375 1.2325 ;
      RECT 64.305 1.1325 64.56 1.2025 ;
      RECT 64.305 0.2725 64.375 0.4075 ;
      RECT 64.305 0.3075 64.56 0.3775 ;
      RECT 62.875 0.2725 62.945 1.2325 ;
      RECT 62.23 0.2725 62.3 0.4075 ;
      RECT 62.23 0.3075 62.945 0.3775 ;
      RECT 61.7675 0.2725 61.8375 1.2325 ;
      RECT 62.6 0.6225 62.67 0.7575 ;
      RECT 61.7675 0.665 62.67 0.735 ;
      RECT 61.5825 1.315 62.145 1.385 ;
      RECT 62.075 0.84 62.145 1.385 ;
      RECT 61.5825 0.2725 61.6525 1.385 ;
      RECT 61.3975 1.0975 61.4675 1.2325 ;
      RECT 61.3975 1.1325 61.6525 1.2025 ;
      RECT 61.3975 0.2725 61.4675 0.4075 ;
      RECT 61.3975 0.3075 61.6525 0.3775 ;
      RECT 59.9675 0.2725 60.0375 1.2325 ;
      RECT 59.3225 0.2725 59.3925 0.4075 ;
      RECT 59.3225 0.3075 60.0375 0.3775 ;
      RECT 58.86 0.2725 58.93 1.2325 ;
      RECT 59.6925 0.6225 59.7625 0.7575 ;
      RECT 58.86 0.665 59.7625 0.735 ;
      RECT 58.675 1.315 59.2375 1.385 ;
      RECT 59.1675 0.84 59.2375 1.385 ;
      RECT 58.675 0.2725 58.745 1.385 ;
      RECT 58.49 1.0975 58.56 1.2325 ;
      RECT 58.49 1.1325 58.745 1.2025 ;
      RECT 58.49 0.2725 58.56 0.4075 ;
      RECT 58.49 0.3075 58.745 0.3775 ;
      RECT 57.06 0.2725 57.13 1.2325 ;
      RECT 56.415 0.2725 56.485 0.4075 ;
      RECT 56.415 0.3075 57.13 0.3775 ;
      RECT 55.9525 0.2725 56.0225 1.2325 ;
      RECT 56.785 0.6225 56.855 0.7575 ;
      RECT 55.9525 0.665 56.855 0.735 ;
      RECT 55.7675 1.315 56.33 1.385 ;
      RECT 56.26 0.84 56.33 1.385 ;
      RECT 55.7675 0.2725 55.8375 1.385 ;
      RECT 55.5825 1.0975 55.6525 1.2325 ;
      RECT 55.5825 1.1325 55.8375 1.2025 ;
      RECT 55.5825 0.2725 55.6525 0.4075 ;
      RECT 55.5825 0.3075 55.8375 0.3775 ;
      RECT 54.1525 0.2725 54.2225 1.2325 ;
      RECT 53.5075 0.2725 53.5775 0.4075 ;
      RECT 53.5075 0.3075 54.2225 0.3775 ;
      RECT 53.045 0.2725 53.115 1.2325 ;
      RECT 53.8775 0.6225 53.9475 0.7575 ;
      RECT 53.045 0.665 53.9475 0.735 ;
      RECT 52.86 1.315 53.4225 1.385 ;
      RECT 53.3525 0.84 53.4225 1.385 ;
      RECT 52.86 0.2725 52.93 1.385 ;
      RECT 52.675 1.0975 52.745 1.2325 ;
      RECT 52.675 1.1325 52.93 1.2025 ;
      RECT 52.675 0.2725 52.745 0.4075 ;
      RECT 52.675 0.3075 52.93 0.3775 ;
      RECT 51.245 0.2725 51.315 1.2325 ;
      RECT 50.6 0.2725 50.67 0.4075 ;
      RECT 50.6 0.3075 51.315 0.3775 ;
      RECT 50.1375 0.2725 50.2075 1.2325 ;
      RECT 50.97 0.6225 51.04 0.7575 ;
      RECT 50.1375 0.665 51.04 0.735 ;
      RECT 49.9525 1.315 50.515 1.385 ;
      RECT 50.445 0.84 50.515 1.385 ;
      RECT 49.9525 0.2725 50.0225 1.385 ;
      RECT 49.7675 1.0975 49.8375 1.2325 ;
      RECT 49.7675 1.1325 50.0225 1.2025 ;
      RECT 49.7675 0.2725 49.8375 0.4075 ;
      RECT 49.7675 0.3075 50.0225 0.3775 ;
      RECT 48.3375 0.2725 48.4075 1.2325 ;
      RECT 47.6925 0.2725 47.7625 0.4075 ;
      RECT 47.6925 0.3075 48.4075 0.3775 ;
      RECT 47.23 0.2725 47.3 1.2325 ;
      RECT 48.0625 0.6225 48.1325 0.7575 ;
      RECT 47.23 0.665 48.1325 0.735 ;
      RECT 47.045 1.315 47.6075 1.385 ;
      RECT 47.5375 0.84 47.6075 1.385 ;
      RECT 47.045 0.2725 47.115 1.385 ;
      RECT 46.86 1.0975 46.93 1.2325 ;
      RECT 46.86 1.1325 47.115 1.2025 ;
      RECT 46.86 0.2725 46.93 0.4075 ;
      RECT 46.86 0.3075 47.115 0.3775 ;
      RECT 45.43 0.2725 45.5 1.2325 ;
      RECT 44.785 0.2725 44.855 0.4075 ;
      RECT 44.785 0.3075 45.5 0.3775 ;
      RECT 44.3225 0.2725 44.3925 1.2325 ;
      RECT 45.155 0.6225 45.225 0.7575 ;
      RECT 44.3225 0.665 45.225 0.735 ;
      RECT 44.1375 1.315 44.7 1.385 ;
      RECT 44.63 0.84 44.7 1.385 ;
      RECT 44.1375 0.2725 44.2075 1.385 ;
      RECT 43.9525 1.0975 44.0225 1.2325 ;
      RECT 43.9525 1.1325 44.2075 1.2025 ;
      RECT 43.9525 0.2725 44.0225 0.4075 ;
      RECT 43.9525 0.3075 44.2075 0.3775 ;
      RECT 42.5225 0.2725 42.5925 1.2325 ;
      RECT 41.8775 0.2725 41.9475 0.4075 ;
      RECT 41.8775 0.3075 42.5925 0.3775 ;
      RECT 41.415 0.2725 41.485 1.2325 ;
      RECT 42.2475 0.6225 42.3175 0.7575 ;
      RECT 41.415 0.665 42.3175 0.735 ;
      RECT 41.23 1.315 41.7925 1.385 ;
      RECT 41.7225 0.84 41.7925 1.385 ;
      RECT 41.23 0.2725 41.3 1.385 ;
      RECT 41.045 1.0975 41.115 1.2325 ;
      RECT 41.045 1.1325 41.3 1.2025 ;
      RECT 41.045 0.2725 41.115 0.4075 ;
      RECT 41.045 0.3075 41.3 0.3775 ;
      RECT 39.615 0.2725 39.685 1.2325 ;
      RECT 38.97 0.2725 39.04 0.4075 ;
      RECT 38.97 0.3075 39.685 0.3775 ;
      RECT 38.5075 0.2725 38.5775 1.2325 ;
      RECT 39.34 0.6225 39.41 0.7575 ;
      RECT 38.5075 0.665 39.41 0.735 ;
      RECT 38.3225 1.315 38.885 1.385 ;
      RECT 38.815 0.84 38.885 1.385 ;
      RECT 38.3225 0.2725 38.3925 1.385 ;
      RECT 38.1375 1.0975 38.2075 1.2325 ;
      RECT 38.1375 1.1325 38.3925 1.2025 ;
      RECT 38.1375 0.2725 38.2075 0.4075 ;
      RECT 38.1375 0.3075 38.3925 0.3775 ;
      RECT 36.7075 0.2725 36.7775 1.2325 ;
      RECT 36.0625 0.2725 36.1325 0.4075 ;
      RECT 36.0625 0.3075 36.7775 0.3775 ;
      RECT 35.6 0.2725 35.67 1.2325 ;
      RECT 36.4325 0.6225 36.5025 0.7575 ;
      RECT 35.6 0.665 36.5025 0.735 ;
      RECT 35.415 1.315 35.9775 1.385 ;
      RECT 35.9075 0.84 35.9775 1.385 ;
      RECT 35.415 0.2725 35.485 1.385 ;
      RECT 35.23 1.0975 35.3 1.2325 ;
      RECT 35.23 1.1325 35.485 1.2025 ;
      RECT 35.23 0.2725 35.3 0.4075 ;
      RECT 35.23 0.3075 35.485 0.3775 ;
      RECT 33.8 0.2725 33.87 1.2325 ;
      RECT 33.155 0.2725 33.225 0.4075 ;
      RECT 33.155 0.3075 33.87 0.3775 ;
      RECT 32.6925 0.2725 32.7625 1.2325 ;
      RECT 33.525 0.6225 33.595 0.7575 ;
      RECT 32.6925 0.665 33.595 0.735 ;
      RECT 32.5075 1.315 33.07 1.385 ;
      RECT 33 0.84 33.07 1.385 ;
      RECT 32.5075 0.2725 32.5775 1.385 ;
      RECT 32.3225 1.0975 32.3925 1.2325 ;
      RECT 32.3225 1.1325 32.5775 1.2025 ;
      RECT 32.3225 0.2725 32.3925 0.4075 ;
      RECT 32.3225 0.3075 32.5775 0.3775 ;
      RECT 30.8925 0.2725 30.9625 1.2325 ;
      RECT 30.2475 0.2725 30.3175 0.4075 ;
      RECT 30.2475 0.3075 30.9625 0.3775 ;
      RECT 29.785 0.2725 29.855 1.2325 ;
      RECT 30.6175 0.6225 30.6875 0.7575 ;
      RECT 29.785 0.665 30.6875 0.735 ;
      RECT 29.6 1.315 30.1625 1.385 ;
      RECT 30.0925 0.84 30.1625 1.385 ;
      RECT 29.6 0.2725 29.67 1.385 ;
      RECT 29.415 1.0975 29.485 1.2325 ;
      RECT 29.415 1.1325 29.67 1.2025 ;
      RECT 29.415 0.2725 29.485 0.4075 ;
      RECT 29.415 0.3075 29.67 0.3775 ;
      RECT 27.985 0.2725 28.055 1.2325 ;
      RECT 27.34 0.2725 27.41 0.4075 ;
      RECT 27.34 0.3075 28.055 0.3775 ;
      RECT 26.8775 0.2725 26.9475 1.2325 ;
      RECT 27.71 0.6225 27.78 0.7575 ;
      RECT 26.8775 0.665 27.78 0.735 ;
      RECT 26.6925 1.315 27.255 1.385 ;
      RECT 27.185 0.84 27.255 1.385 ;
      RECT 26.6925 0.2725 26.7625 1.385 ;
      RECT 26.5075 1.0975 26.5775 1.2325 ;
      RECT 26.5075 1.1325 26.7625 1.2025 ;
      RECT 26.5075 0.2725 26.5775 0.4075 ;
      RECT 26.5075 0.3075 26.7625 0.3775 ;
      RECT 25.0775 0.2725 25.1475 1.2325 ;
      RECT 24.4325 0.2725 24.5025 0.4075 ;
      RECT 24.4325 0.3075 25.1475 0.3775 ;
      RECT 23.97 0.2725 24.04 1.2325 ;
      RECT 24.8025 0.6225 24.8725 0.7575 ;
      RECT 23.97 0.665 24.8725 0.735 ;
      RECT 23.785 1.315 24.3475 1.385 ;
      RECT 24.2775 0.84 24.3475 1.385 ;
      RECT 23.785 0.2725 23.855 1.385 ;
      RECT 23.6 1.0975 23.67 1.2325 ;
      RECT 23.6 1.1325 23.855 1.2025 ;
      RECT 23.6 0.2725 23.67 0.4075 ;
      RECT 23.6 0.3075 23.855 0.3775 ;
      RECT 22.17 0.2725 22.24 1.2325 ;
      RECT 21.525 0.2725 21.595 0.4075 ;
      RECT 21.525 0.3075 22.24 0.3775 ;
      RECT 21.0625 0.2725 21.1325 1.2325 ;
      RECT 21.895 0.6225 21.965 0.7575 ;
      RECT 21.0625 0.665 21.965 0.735 ;
      RECT 20.8775 1.315 21.44 1.385 ;
      RECT 21.37 0.84 21.44 1.385 ;
      RECT 20.8775 0.2725 20.9475 1.385 ;
      RECT 20.6925 1.0975 20.7625 1.2325 ;
      RECT 20.6925 1.1325 20.9475 1.2025 ;
      RECT 20.6925 0.2725 20.7625 0.4075 ;
      RECT 20.6925 0.3075 20.9475 0.3775 ;
      RECT 19.2625 0.2725 19.3325 1.2325 ;
      RECT 18.6175 0.2725 18.6875 0.4075 ;
      RECT 18.6175 0.3075 19.3325 0.3775 ;
      RECT 18.155 0.2725 18.225 1.2325 ;
      RECT 18.9875 0.6225 19.0575 0.7575 ;
      RECT 18.155 0.665 19.0575 0.735 ;
      RECT 17.97 1.315 18.5325 1.385 ;
      RECT 18.4625 0.84 18.5325 1.385 ;
      RECT 17.97 0.2725 18.04 1.385 ;
      RECT 17.785 1.0975 17.855 1.2325 ;
      RECT 17.785 1.1325 18.04 1.2025 ;
      RECT 17.785 0.2725 17.855 0.4075 ;
      RECT 17.785 0.3075 18.04 0.3775 ;
      RECT 16.355 0.2725 16.425 1.2325 ;
      RECT 15.71 0.2725 15.78 0.4075 ;
      RECT 15.71 0.3075 16.425 0.3775 ;
      RECT 15.2475 0.2725 15.3175 1.2325 ;
      RECT 16.08 0.6225 16.15 0.7575 ;
      RECT 15.2475 0.665 16.15 0.735 ;
      RECT 15.0625 1.315 15.625 1.385 ;
      RECT 15.555 0.84 15.625 1.385 ;
      RECT 15.0625 0.2725 15.1325 1.385 ;
      RECT 14.8775 1.0975 14.9475 1.2325 ;
      RECT 14.8775 1.1325 15.1325 1.2025 ;
      RECT 14.8775 0.2725 14.9475 0.4075 ;
      RECT 14.8775 0.3075 15.1325 0.3775 ;
      RECT 13.4475 0.2725 13.5175 1.2325 ;
      RECT 12.8025 0.2725 12.8725 0.4075 ;
      RECT 12.8025 0.3075 13.5175 0.3775 ;
      RECT 12.34 0.2725 12.41 1.2325 ;
      RECT 13.1725 0.6225 13.2425 0.7575 ;
      RECT 12.34 0.665 13.2425 0.735 ;
      RECT 12.155 1.315 12.7175 1.385 ;
      RECT 12.6475 0.84 12.7175 1.385 ;
      RECT 12.155 0.2725 12.225 1.385 ;
      RECT 11.97 1.0975 12.04 1.2325 ;
      RECT 11.97 1.1325 12.225 1.2025 ;
      RECT 11.97 0.2725 12.04 0.4075 ;
      RECT 11.97 0.3075 12.225 0.3775 ;
      RECT 10.54 0.2725 10.61 1.2325 ;
      RECT 9.895 0.2725 9.965 0.4075 ;
      RECT 9.895 0.3075 10.61 0.3775 ;
      RECT 9.4325 0.2725 9.5025 1.2325 ;
      RECT 10.265 0.6225 10.335 0.7575 ;
      RECT 9.4325 0.665 10.335 0.735 ;
      RECT 9.2475 1.315 9.81 1.385 ;
      RECT 9.74 0.84 9.81 1.385 ;
      RECT 9.2475 0.2725 9.3175 1.385 ;
      RECT 9.0625 1.0975 9.1325 1.2325 ;
      RECT 9.0625 1.1325 9.3175 1.2025 ;
      RECT 9.0625 0.2725 9.1325 0.4075 ;
      RECT 9.0625 0.3075 9.3175 0.3775 ;
      RECT 7.6325 0.2725 7.7025 1.2325 ;
      RECT 6.9875 0.2725 7.0575 0.4075 ;
      RECT 6.9875 0.3075 7.7025 0.3775 ;
      RECT 6.525 0.2725 6.595 1.2325 ;
      RECT 7.3575 0.6225 7.4275 0.7575 ;
      RECT 6.525 0.665 7.4275 0.735 ;
      RECT 6.34 1.315 6.9025 1.385 ;
      RECT 6.8325 0.84 6.9025 1.385 ;
      RECT 6.34 0.2725 6.41 1.385 ;
      RECT 6.155 1.0975 6.225 1.2325 ;
      RECT 6.155 1.1325 6.41 1.2025 ;
      RECT 6.155 0.2725 6.225 0.4075 ;
      RECT 6.155 0.3075 6.41 0.3775 ;
      RECT 4.725 0.2725 4.795 1.2325 ;
      RECT 4.08 0.2725 4.15 0.4075 ;
      RECT 4.08 0.3075 4.795 0.3775 ;
      RECT 3.6175 0.2725 3.6875 1.2325 ;
      RECT 4.45 0.6225 4.52 0.7575 ;
      RECT 3.6175 0.665 4.52 0.735 ;
      RECT 3.4325 1.315 3.995 1.385 ;
      RECT 3.925 0.84 3.995 1.385 ;
      RECT 3.4325 0.2725 3.5025 1.385 ;
      RECT 3.2475 1.0975 3.3175 1.2325 ;
      RECT 3.2475 1.1325 3.5025 1.2025 ;
      RECT 3.2475 0.2725 3.3175 0.4075 ;
      RECT 3.2475 0.3075 3.5025 0.3775 ;
      RECT 1.8175 0.2725 1.8875 1.2325 ;
      RECT 1.1725 0.2725 1.2425 0.4075 ;
      RECT 1.1725 0.3075 1.8875 0.3775 ;
      RECT 0.71 0.2725 0.78 1.2325 ;
      RECT 1.5425 0.6225 1.6125 0.7575 ;
      RECT 0.71 0.665 1.6125 0.735 ;
      RECT 0.525 1.315 1.0875 1.385 ;
      RECT 1.0175 0.84 1.0875 1.385 ;
      RECT 0.525 0.2725 0.595 1.385 ;
      RECT 0.34 1.0975 0.41 1.2325 ;
      RECT 0.34 1.1325 0.595 1.2025 ;
      RECT 0.34 0.2725 0.41 0.4075 ;
      RECT 0.34 0.3075 0.595 0.3775 ;
      RECT 95.295 0.2725 95.365 1.2325 ;
      RECT 94.9125 0.2675 94.9825 1.2325 ;
      RECT 93.8575 0.75 93.9275 0.89 ;
      RECT 93.265 0.2725 93.335 1.2325 ;
      RECT 92.8825 0.2675 92.9525 1.2325 ;
      RECT 91.8275 0.75 91.8975 0.89 ;
      RECT 91.4925 0.2725 91.5625 1.235 ;
      RECT 91.3075 0.2725 91.3775 1.2325 ;
      RECT 90.835 0.27 90.905 1.2325 ;
      RECT 90.65 0.2725 90.72 1.2325 ;
      RECT 89.885 0.2725 89.955 1.235 ;
      RECT 89.7 0.2725 89.77 1.2325 ;
      RECT 89.2275 0.27 89.2975 1.2325 ;
      RECT 86.9775 0.2725 87.0475 1.235 ;
      RECT 86.7925 0.2725 86.8625 1.2325 ;
      RECT 86.32 0.27 86.39 1.2325 ;
      RECT 84.07 0.2725 84.14 1.235 ;
      RECT 83.885 0.2725 83.955 1.2325 ;
      RECT 83.4125 0.27 83.4825 1.2325 ;
      RECT 81.1625 0.2725 81.2325 1.235 ;
      RECT 80.9775 0.2725 81.0475 1.2325 ;
      RECT 80.505 0.27 80.575 1.2325 ;
      RECT 78.255 0.2725 78.325 1.235 ;
      RECT 78.07 0.2725 78.14 1.2325 ;
      RECT 77.5975 0.27 77.6675 1.2325 ;
      RECT 75.3475 0.2725 75.4175 1.235 ;
      RECT 75.1625 0.2725 75.2325 1.2325 ;
      RECT 74.69 0.27 74.76 1.2325 ;
      RECT 72.44 0.2725 72.51 1.235 ;
      RECT 72.255 0.2725 72.325 1.2325 ;
      RECT 71.7825 0.27 71.8525 1.2325 ;
      RECT 69.5325 0.2725 69.6025 1.235 ;
      RECT 69.3475 0.2725 69.4175 1.2325 ;
      RECT 68.875 0.27 68.945 1.2325 ;
      RECT 66.625 0.2725 66.695 1.235 ;
      RECT 66.44 0.2725 66.51 1.2325 ;
      RECT 65.9675 0.27 66.0375 1.2325 ;
      RECT 63.7175 0.2725 63.7875 1.235 ;
      RECT 63.5325 0.2725 63.6025 1.2325 ;
      RECT 63.06 0.27 63.13 1.2325 ;
      RECT 60.81 0.2725 60.88 1.235 ;
      RECT 60.625 0.2725 60.695 1.2325 ;
      RECT 60.1525 0.27 60.2225 1.2325 ;
      RECT 57.9025 0.2725 57.9725 1.235 ;
      RECT 57.7175 0.2725 57.7875 1.2325 ;
      RECT 57.245 0.27 57.315 1.2325 ;
      RECT 54.995 0.2725 55.065 1.235 ;
      RECT 54.81 0.2725 54.88 1.2325 ;
      RECT 54.3375 0.27 54.4075 1.2325 ;
      RECT 52.0875 0.2725 52.1575 1.235 ;
      RECT 51.9025 0.2725 51.9725 1.2325 ;
      RECT 51.43 0.27 51.5 1.2325 ;
      RECT 49.18 0.2725 49.25 1.235 ;
      RECT 48.995 0.2725 49.065 1.2325 ;
      RECT 48.5225 0.27 48.5925 1.2325 ;
      RECT 46.2725 0.2725 46.3425 1.235 ;
      RECT 46.0875 0.2725 46.1575 1.2325 ;
      RECT 45.615 0.27 45.685 1.2325 ;
      RECT 43.365 0.2725 43.435 1.235 ;
      RECT 43.18 0.2725 43.25 1.2325 ;
      RECT 42.7075 0.27 42.7775 1.2325 ;
      RECT 40.4575 0.2725 40.5275 1.235 ;
      RECT 40.2725 0.2725 40.3425 1.2325 ;
      RECT 39.8 0.27 39.87 1.2325 ;
      RECT 37.55 0.2725 37.62 1.235 ;
      RECT 37.365 0.2725 37.435 1.2325 ;
      RECT 36.8925 0.27 36.9625 1.2325 ;
      RECT 34.6425 0.2725 34.7125 1.235 ;
      RECT 34.4575 0.2725 34.5275 1.2325 ;
      RECT 33.985 0.27 34.055 1.2325 ;
      RECT 31.735 0.2725 31.805 1.235 ;
      RECT 31.55 0.2725 31.62 1.2325 ;
      RECT 31.0775 0.27 31.1475 1.2325 ;
      RECT 28.8275 0.2725 28.8975 1.235 ;
      RECT 28.6425 0.2725 28.7125 1.2325 ;
      RECT 28.17 0.27 28.24 1.2325 ;
      RECT 25.92 0.2725 25.99 1.235 ;
      RECT 25.735 0.2725 25.805 1.2325 ;
      RECT 25.2625 0.27 25.3325 1.2325 ;
      RECT 23.0125 0.2725 23.0825 1.235 ;
      RECT 22.8275 0.2725 22.8975 1.2325 ;
      RECT 22.355 0.27 22.425 1.2325 ;
      RECT 20.105 0.2725 20.175 1.235 ;
      RECT 19.92 0.2725 19.99 1.2325 ;
      RECT 19.4475 0.27 19.5175 1.2325 ;
      RECT 17.1975 0.2725 17.2675 1.235 ;
      RECT 17.0125 0.2725 17.0825 1.2325 ;
      RECT 16.54 0.27 16.61 1.2325 ;
      RECT 14.29 0.2725 14.36 1.235 ;
      RECT 14.105 0.2725 14.175 1.2325 ;
      RECT 13.6325 0.27 13.7025 1.2325 ;
      RECT 11.3825 0.2725 11.4525 1.235 ;
      RECT 11.1975 0.2725 11.2675 1.2325 ;
      RECT 10.725 0.27 10.795 1.2325 ;
      RECT 8.475 0.2725 8.545 1.235 ;
      RECT 8.29 0.2725 8.36 1.2325 ;
      RECT 7.8175 0.27 7.8875 1.2325 ;
      RECT 5.5675 0.2725 5.6375 1.235 ;
      RECT 5.3825 0.2725 5.4525 1.2325 ;
      RECT 4.91 0.27 4.98 1.2325 ;
      RECT 2.66 0.2725 2.73 1.235 ;
      RECT 2.475 0.2725 2.545 1.2325 ;
      RECT 2.0025 0.27 2.0725 1.2325 ;
    LAYER metal3 ;
      RECT 93.8575 0.75 93.9275 0.89 ;
      RECT 91.8275 0.75 91.8975 0.89 ;
      RECT 91.4925 1.095 91.5625 1.235 ;
      RECT 90.835 0.27 90.905 0.41 ;
      RECT 89.885 1.095 89.955 1.235 ;
      RECT 89.2275 0.27 89.2975 0.41 ;
      RECT 86.9775 1.095 87.0475 1.235 ;
      RECT 86.32 0.27 86.39 0.41 ;
      RECT 84.07 1.095 84.14 1.235 ;
      RECT 83.4125 0.27 83.4825 0.41 ;
      RECT 81.1625 1.095 81.2325 1.235 ;
      RECT 80.505 0.27 80.575 0.41 ;
      RECT 78.255 1.095 78.325 1.235 ;
      RECT 77.5975 0.27 77.6675 0.41 ;
      RECT 75.3475 1.095 75.4175 1.235 ;
      RECT 74.69 0.27 74.76 0.41 ;
      RECT 72.44 1.095 72.51 1.235 ;
      RECT 71.7825 0.27 71.8525 0.41 ;
      RECT 69.5325 1.095 69.6025 1.235 ;
      RECT 68.875 0.27 68.945 0.41 ;
      RECT 66.625 1.095 66.695 1.235 ;
      RECT 65.9675 0.27 66.0375 0.41 ;
      RECT 63.7175 1.095 63.7875 1.235 ;
      RECT 63.06 0.27 63.13 0.41 ;
      RECT 60.81 1.095 60.88 1.235 ;
      RECT 60.1525 0.27 60.2225 0.41 ;
      RECT 57.9025 1.095 57.9725 1.235 ;
      RECT 57.245 0.27 57.315 0.41 ;
      RECT 54.995 1.095 55.065 1.235 ;
      RECT 54.3375 0.27 54.4075 0.41 ;
      RECT 52.0875 1.095 52.1575 1.235 ;
      RECT 51.43 0.27 51.5 0.41 ;
      RECT 49.18 1.095 49.25 1.235 ;
      RECT 48.5225 0.27 48.5925 0.41 ;
      RECT 46.2725 1.095 46.3425 1.235 ;
      RECT 45.615 0.27 45.685 0.41 ;
      RECT 43.365 1.095 43.435 1.235 ;
      RECT 42.7075 0.27 42.7775 0.41 ;
      RECT 40.4575 1.095 40.5275 1.235 ;
      RECT 39.8 0.27 39.87 0.41 ;
      RECT 37.55 1.095 37.62 1.235 ;
      RECT 36.8925 0.27 36.9625 0.41 ;
      RECT 34.6425 1.095 34.7125 1.235 ;
      RECT 33.985 0.27 34.055 0.41 ;
      RECT 31.735 1.095 31.805 1.235 ;
      RECT 31.0775 0.27 31.1475 0.41 ;
      RECT 28.8275 1.095 28.8975 1.235 ;
      RECT 28.17 0.27 28.24 0.41 ;
      RECT 25.92 1.095 25.99 1.235 ;
      RECT 25.2625 0.27 25.3325 0.41 ;
      RECT 23.0125 1.095 23.0825 1.235 ;
      RECT 22.355 0.27 22.425 0.41 ;
      RECT 20.105 1.095 20.175 1.235 ;
      RECT 19.4475 0.27 19.5175 0.41 ;
      RECT 17.1975 1.095 17.2675 1.235 ;
      RECT 16.54 0.27 16.61 0.41 ;
      RECT 14.29 1.095 14.36 1.235 ;
      RECT 13.6325 0.27 13.7025 0.41 ;
      RECT 11.3825 1.095 11.4525 1.235 ;
      RECT 10.725 0.27 10.795 0.41 ;
      RECT 8.475 1.095 8.545 1.235 ;
      RECT 7.8175 0.27 7.8875 0.41 ;
      RECT 5.5675 1.095 5.6375 1.235 ;
      RECT 4.91 0.27 4.98 0.41 ;
      RECT 2.66 1.095 2.73 1.235 ;
      RECT 2.0025 0.27 2.0725 0.41 ;
    LAYER metal4 ;
      RECT 93.8225 0.75 93.965 0.89 ;
      RECT 93.825 0.27 93.965 0.89 ;
      RECT 1.9675 0.27 93.965 0.41 ;
      RECT 2.625 1.095 91.9325 1.235 ;
      RECT 91.7925 0.75 91.9325 1.235 ;
    LAYER via1 ;
      RECT 95.535 0.82 95.6 0.885 ;
      RECT 95.2975 0.3075 95.3625 0.3725 ;
      RECT 95.2975 1.1325 95.3625 1.1975 ;
      RECT 95.105 0.3075 95.17 0.3725 ;
      RECT 95.105 1.1325 95.17 1.1975 ;
      RECT 94.915 0.3075 94.98 0.3725 ;
      RECT 94.915 1.1325 94.98 1.1975 ;
      RECT 94.715 0.7425 94.78 0.8075 ;
      RECT 94.0175 0.525 94.0825 0.59 ;
      RECT 93.86 0.7875 93.925 0.8525 ;
      RECT 93.505 0.82 93.57 0.885 ;
      RECT 93.2675 0.3075 93.3325 0.3725 ;
      RECT 93.2675 1.1325 93.3325 1.1975 ;
      RECT 93.075 0.3075 93.14 0.3725 ;
      RECT 93.075 1.1325 93.14 1.1975 ;
      RECT 92.885 0.3075 92.95 0.3725 ;
      RECT 92.885 1.1325 92.95 1.1975 ;
      RECT 92.685 0.7425 92.75 0.8075 ;
      RECT 91.9875 0.525 92.0525 0.59 ;
      RECT 91.83 0.7875 91.895 0.8525 ;
      RECT 91.495 0.3075 91.56 0.3725 ;
      RECT 91.495 1.1325 91.56 1.1975 ;
      RECT 91.31 0.3075 91.375 0.3725 ;
      RECT 91.31 0.6925 91.375 0.7575 ;
      RECT 91.31 1.1325 91.375 1.1975 ;
      RECT 90.8375 0.3075 90.9025 0.3725 ;
      RECT 90.8375 1.1325 90.9025 1.1975 ;
      RECT 90.6525 0.3075 90.7175 0.3725 ;
      RECT 90.6525 0.6825 90.7175 0.7475 ;
      RECT 90.6525 1.1325 90.7175 1.1975 ;
      RECT 89.8875 0.3075 89.9525 0.3725 ;
      RECT 89.8875 1.1325 89.9525 1.1975 ;
      RECT 89.7025 0.3075 89.7675 0.3725 ;
      RECT 89.7025 0.6925 89.7675 0.7575 ;
      RECT 89.7025 1.1325 89.7675 1.1975 ;
      RECT 89.23 0.3075 89.295 0.3725 ;
      RECT 89.23 1.1325 89.295 1.1975 ;
      RECT 89.045 0.3075 89.11 0.3725 ;
      RECT 89.045 0.6825 89.11 0.7475 ;
      RECT 89.045 1.1325 89.11 1.1975 ;
      RECT 88.77 0.6575 88.835 0.7225 ;
      RECT 88.4 0.3075 88.465 0.3725 ;
      RECT 88.245 0.875 88.31 0.94 ;
      RECT 87.9375 0.3075 88.0025 0.3725 ;
      RECT 87.9375 1.1325 88.0025 1.1975 ;
      RECT 87.7525 0.3075 87.8175 0.3725 ;
      RECT 87.7525 1.1325 87.8175 1.1975 ;
      RECT 87.5675 0.3075 87.6325 0.3725 ;
      RECT 87.5675 1.1325 87.6325 1.1975 ;
      RECT 86.98 0.3075 87.045 0.3725 ;
      RECT 86.98 1.1325 87.045 1.1975 ;
      RECT 86.795 0.3075 86.86 0.3725 ;
      RECT 86.795 0.6925 86.86 0.7575 ;
      RECT 86.795 1.1325 86.86 1.1975 ;
      RECT 86.3225 0.3075 86.3875 0.3725 ;
      RECT 86.3225 1.1325 86.3875 1.1975 ;
      RECT 86.1375 0.3075 86.2025 0.3725 ;
      RECT 86.1375 0.6825 86.2025 0.7475 ;
      RECT 86.1375 1.1325 86.2025 1.1975 ;
      RECT 85.8625 0.6575 85.9275 0.7225 ;
      RECT 85.4925 0.3075 85.5575 0.3725 ;
      RECT 85.3375 0.875 85.4025 0.94 ;
      RECT 85.03 0.3075 85.095 0.3725 ;
      RECT 85.03 1.1325 85.095 1.1975 ;
      RECT 84.845 0.3075 84.91 0.3725 ;
      RECT 84.845 1.1325 84.91 1.1975 ;
      RECT 84.66 0.3075 84.725 0.3725 ;
      RECT 84.66 1.1325 84.725 1.1975 ;
      RECT 84.0725 0.3075 84.1375 0.3725 ;
      RECT 84.0725 1.1325 84.1375 1.1975 ;
      RECT 83.8875 0.3075 83.9525 0.3725 ;
      RECT 83.8875 0.6925 83.9525 0.7575 ;
      RECT 83.8875 1.1325 83.9525 1.1975 ;
      RECT 83.415 0.3075 83.48 0.3725 ;
      RECT 83.415 1.1325 83.48 1.1975 ;
      RECT 83.23 0.3075 83.295 0.3725 ;
      RECT 83.23 0.6825 83.295 0.7475 ;
      RECT 83.23 1.1325 83.295 1.1975 ;
      RECT 82.955 0.6575 83.02 0.7225 ;
      RECT 82.585 0.3075 82.65 0.3725 ;
      RECT 82.43 0.875 82.495 0.94 ;
      RECT 82.1225 0.3075 82.1875 0.3725 ;
      RECT 82.1225 1.1325 82.1875 1.1975 ;
      RECT 81.9375 0.3075 82.0025 0.3725 ;
      RECT 81.9375 1.1325 82.0025 1.1975 ;
      RECT 81.7525 0.3075 81.8175 0.3725 ;
      RECT 81.7525 1.1325 81.8175 1.1975 ;
      RECT 81.165 0.3075 81.23 0.3725 ;
      RECT 81.165 1.1325 81.23 1.1975 ;
      RECT 80.98 0.3075 81.045 0.3725 ;
      RECT 80.98 0.6925 81.045 0.7575 ;
      RECT 80.98 1.1325 81.045 1.1975 ;
      RECT 80.5075 0.3075 80.5725 0.3725 ;
      RECT 80.5075 1.1325 80.5725 1.1975 ;
      RECT 80.3225 0.3075 80.3875 0.3725 ;
      RECT 80.3225 0.6825 80.3875 0.7475 ;
      RECT 80.3225 1.1325 80.3875 1.1975 ;
      RECT 80.0475 0.6575 80.1125 0.7225 ;
      RECT 79.6775 0.3075 79.7425 0.3725 ;
      RECT 79.5225 0.875 79.5875 0.94 ;
      RECT 79.215 0.3075 79.28 0.3725 ;
      RECT 79.215 1.1325 79.28 1.1975 ;
      RECT 79.03 0.3075 79.095 0.3725 ;
      RECT 79.03 1.1325 79.095 1.1975 ;
      RECT 78.845 0.3075 78.91 0.3725 ;
      RECT 78.845 1.1325 78.91 1.1975 ;
      RECT 78.2575 0.3075 78.3225 0.3725 ;
      RECT 78.2575 1.1325 78.3225 1.1975 ;
      RECT 78.0725 0.3075 78.1375 0.3725 ;
      RECT 78.0725 0.6925 78.1375 0.7575 ;
      RECT 78.0725 1.1325 78.1375 1.1975 ;
      RECT 77.6 0.3075 77.665 0.3725 ;
      RECT 77.6 1.1325 77.665 1.1975 ;
      RECT 77.415 0.3075 77.48 0.3725 ;
      RECT 77.415 0.6825 77.48 0.7475 ;
      RECT 77.415 1.1325 77.48 1.1975 ;
      RECT 77.14 0.6575 77.205 0.7225 ;
      RECT 76.77 0.3075 76.835 0.3725 ;
      RECT 76.615 0.875 76.68 0.94 ;
      RECT 76.3075 0.3075 76.3725 0.3725 ;
      RECT 76.3075 1.1325 76.3725 1.1975 ;
      RECT 76.1225 0.3075 76.1875 0.3725 ;
      RECT 76.1225 1.1325 76.1875 1.1975 ;
      RECT 75.9375 0.3075 76.0025 0.3725 ;
      RECT 75.9375 1.1325 76.0025 1.1975 ;
      RECT 75.35 0.3075 75.415 0.3725 ;
      RECT 75.35 1.1325 75.415 1.1975 ;
      RECT 75.165 0.3075 75.23 0.3725 ;
      RECT 75.165 0.6925 75.23 0.7575 ;
      RECT 75.165 1.1325 75.23 1.1975 ;
      RECT 74.6925 0.3075 74.7575 0.3725 ;
      RECT 74.6925 1.1325 74.7575 1.1975 ;
      RECT 74.5075 0.3075 74.5725 0.3725 ;
      RECT 74.5075 0.6825 74.5725 0.7475 ;
      RECT 74.5075 1.1325 74.5725 1.1975 ;
      RECT 74.2325 0.6575 74.2975 0.7225 ;
      RECT 73.8625 0.3075 73.9275 0.3725 ;
      RECT 73.7075 0.875 73.7725 0.94 ;
      RECT 73.4 0.3075 73.465 0.3725 ;
      RECT 73.4 1.1325 73.465 1.1975 ;
      RECT 73.215 0.3075 73.28 0.3725 ;
      RECT 73.215 1.1325 73.28 1.1975 ;
      RECT 73.03 0.3075 73.095 0.3725 ;
      RECT 73.03 1.1325 73.095 1.1975 ;
      RECT 72.4425 0.3075 72.5075 0.3725 ;
      RECT 72.4425 1.1325 72.5075 1.1975 ;
      RECT 72.2575 0.3075 72.3225 0.3725 ;
      RECT 72.2575 0.6925 72.3225 0.7575 ;
      RECT 72.2575 1.1325 72.3225 1.1975 ;
      RECT 71.785 0.3075 71.85 0.3725 ;
      RECT 71.785 1.1325 71.85 1.1975 ;
      RECT 71.6 0.3075 71.665 0.3725 ;
      RECT 71.6 0.6825 71.665 0.7475 ;
      RECT 71.6 1.1325 71.665 1.1975 ;
      RECT 71.325 0.6575 71.39 0.7225 ;
      RECT 70.955 0.3075 71.02 0.3725 ;
      RECT 70.8 0.875 70.865 0.94 ;
      RECT 70.4925 0.3075 70.5575 0.3725 ;
      RECT 70.4925 1.1325 70.5575 1.1975 ;
      RECT 70.3075 0.3075 70.3725 0.3725 ;
      RECT 70.3075 1.1325 70.3725 1.1975 ;
      RECT 70.1225 0.3075 70.1875 0.3725 ;
      RECT 70.1225 1.1325 70.1875 1.1975 ;
      RECT 69.535 0.3075 69.6 0.3725 ;
      RECT 69.535 1.1325 69.6 1.1975 ;
      RECT 69.35 0.3075 69.415 0.3725 ;
      RECT 69.35 0.6925 69.415 0.7575 ;
      RECT 69.35 1.1325 69.415 1.1975 ;
      RECT 68.8775 0.3075 68.9425 0.3725 ;
      RECT 68.8775 1.1325 68.9425 1.1975 ;
      RECT 68.6925 0.3075 68.7575 0.3725 ;
      RECT 68.6925 0.6825 68.7575 0.7475 ;
      RECT 68.6925 1.1325 68.7575 1.1975 ;
      RECT 68.4175 0.6575 68.4825 0.7225 ;
      RECT 68.0475 0.3075 68.1125 0.3725 ;
      RECT 67.8925 0.875 67.9575 0.94 ;
      RECT 67.585 0.3075 67.65 0.3725 ;
      RECT 67.585 1.1325 67.65 1.1975 ;
      RECT 67.4 0.3075 67.465 0.3725 ;
      RECT 67.4 1.1325 67.465 1.1975 ;
      RECT 67.215 0.3075 67.28 0.3725 ;
      RECT 67.215 1.1325 67.28 1.1975 ;
      RECT 66.6275 0.3075 66.6925 0.3725 ;
      RECT 66.6275 1.1325 66.6925 1.1975 ;
      RECT 66.4425 0.3075 66.5075 0.3725 ;
      RECT 66.4425 0.6925 66.5075 0.7575 ;
      RECT 66.4425 1.1325 66.5075 1.1975 ;
      RECT 65.97 0.3075 66.035 0.3725 ;
      RECT 65.97 1.1325 66.035 1.1975 ;
      RECT 65.785 0.3075 65.85 0.3725 ;
      RECT 65.785 0.6825 65.85 0.7475 ;
      RECT 65.785 1.1325 65.85 1.1975 ;
      RECT 65.51 0.6575 65.575 0.7225 ;
      RECT 65.14 0.3075 65.205 0.3725 ;
      RECT 64.985 0.875 65.05 0.94 ;
      RECT 64.6775 0.3075 64.7425 0.3725 ;
      RECT 64.6775 1.1325 64.7425 1.1975 ;
      RECT 64.4925 0.3075 64.5575 0.3725 ;
      RECT 64.4925 1.1325 64.5575 1.1975 ;
      RECT 64.3075 0.3075 64.3725 0.3725 ;
      RECT 64.3075 1.1325 64.3725 1.1975 ;
      RECT 63.72 0.3075 63.785 0.3725 ;
      RECT 63.72 1.1325 63.785 1.1975 ;
      RECT 63.535 0.3075 63.6 0.3725 ;
      RECT 63.535 0.6925 63.6 0.7575 ;
      RECT 63.535 1.1325 63.6 1.1975 ;
      RECT 63.0625 0.3075 63.1275 0.3725 ;
      RECT 63.0625 1.1325 63.1275 1.1975 ;
      RECT 62.8775 0.3075 62.9425 0.3725 ;
      RECT 62.8775 0.6825 62.9425 0.7475 ;
      RECT 62.8775 1.1325 62.9425 1.1975 ;
      RECT 62.6025 0.6575 62.6675 0.7225 ;
      RECT 62.2325 0.3075 62.2975 0.3725 ;
      RECT 62.0775 0.875 62.1425 0.94 ;
      RECT 61.77 0.3075 61.835 0.3725 ;
      RECT 61.77 1.1325 61.835 1.1975 ;
      RECT 61.585 0.3075 61.65 0.3725 ;
      RECT 61.585 1.1325 61.65 1.1975 ;
      RECT 61.4 0.3075 61.465 0.3725 ;
      RECT 61.4 1.1325 61.465 1.1975 ;
      RECT 60.8125 0.3075 60.8775 0.3725 ;
      RECT 60.8125 1.1325 60.8775 1.1975 ;
      RECT 60.6275 0.3075 60.6925 0.3725 ;
      RECT 60.6275 0.6925 60.6925 0.7575 ;
      RECT 60.6275 1.1325 60.6925 1.1975 ;
      RECT 60.155 0.3075 60.22 0.3725 ;
      RECT 60.155 1.1325 60.22 1.1975 ;
      RECT 59.97 0.3075 60.035 0.3725 ;
      RECT 59.97 0.6825 60.035 0.7475 ;
      RECT 59.97 1.1325 60.035 1.1975 ;
      RECT 59.695 0.6575 59.76 0.7225 ;
      RECT 59.325 0.3075 59.39 0.3725 ;
      RECT 59.17 0.875 59.235 0.94 ;
      RECT 58.8625 0.3075 58.9275 0.3725 ;
      RECT 58.8625 1.1325 58.9275 1.1975 ;
      RECT 58.6775 0.3075 58.7425 0.3725 ;
      RECT 58.6775 1.1325 58.7425 1.1975 ;
      RECT 58.4925 0.3075 58.5575 0.3725 ;
      RECT 58.4925 1.1325 58.5575 1.1975 ;
      RECT 57.905 0.3075 57.97 0.3725 ;
      RECT 57.905 1.1325 57.97 1.1975 ;
      RECT 57.72 0.3075 57.785 0.3725 ;
      RECT 57.72 0.6925 57.785 0.7575 ;
      RECT 57.72 1.1325 57.785 1.1975 ;
      RECT 57.2475 0.3075 57.3125 0.3725 ;
      RECT 57.2475 1.1325 57.3125 1.1975 ;
      RECT 57.0625 0.3075 57.1275 0.3725 ;
      RECT 57.0625 0.6825 57.1275 0.7475 ;
      RECT 57.0625 1.1325 57.1275 1.1975 ;
      RECT 56.7875 0.6575 56.8525 0.7225 ;
      RECT 56.4175 0.3075 56.4825 0.3725 ;
      RECT 56.2625 0.875 56.3275 0.94 ;
      RECT 55.955 0.3075 56.02 0.3725 ;
      RECT 55.955 1.1325 56.02 1.1975 ;
      RECT 55.77 0.3075 55.835 0.3725 ;
      RECT 55.77 1.1325 55.835 1.1975 ;
      RECT 55.585 0.3075 55.65 0.3725 ;
      RECT 55.585 1.1325 55.65 1.1975 ;
      RECT 54.9975 0.3075 55.0625 0.3725 ;
      RECT 54.9975 1.1325 55.0625 1.1975 ;
      RECT 54.8125 0.3075 54.8775 0.3725 ;
      RECT 54.8125 0.6925 54.8775 0.7575 ;
      RECT 54.8125 1.1325 54.8775 1.1975 ;
      RECT 54.34 0.3075 54.405 0.3725 ;
      RECT 54.34 1.1325 54.405 1.1975 ;
      RECT 54.155 0.3075 54.22 0.3725 ;
      RECT 54.155 0.6825 54.22 0.7475 ;
      RECT 54.155 1.1325 54.22 1.1975 ;
      RECT 53.88 0.6575 53.945 0.7225 ;
      RECT 53.51 0.3075 53.575 0.3725 ;
      RECT 53.355 0.875 53.42 0.94 ;
      RECT 53.0475 0.3075 53.1125 0.3725 ;
      RECT 53.0475 1.1325 53.1125 1.1975 ;
      RECT 52.8625 0.3075 52.9275 0.3725 ;
      RECT 52.8625 1.1325 52.9275 1.1975 ;
      RECT 52.6775 0.3075 52.7425 0.3725 ;
      RECT 52.6775 1.1325 52.7425 1.1975 ;
      RECT 52.09 0.3075 52.155 0.3725 ;
      RECT 52.09 1.1325 52.155 1.1975 ;
      RECT 51.905 0.3075 51.97 0.3725 ;
      RECT 51.905 0.6925 51.97 0.7575 ;
      RECT 51.905 1.1325 51.97 1.1975 ;
      RECT 51.4325 0.3075 51.4975 0.3725 ;
      RECT 51.4325 1.1325 51.4975 1.1975 ;
      RECT 51.2475 0.3075 51.3125 0.3725 ;
      RECT 51.2475 0.6825 51.3125 0.7475 ;
      RECT 51.2475 1.1325 51.3125 1.1975 ;
      RECT 50.9725 0.6575 51.0375 0.7225 ;
      RECT 50.6025 0.3075 50.6675 0.3725 ;
      RECT 50.4475 0.875 50.5125 0.94 ;
      RECT 50.14 0.3075 50.205 0.3725 ;
      RECT 50.14 1.1325 50.205 1.1975 ;
      RECT 49.955 0.3075 50.02 0.3725 ;
      RECT 49.955 1.1325 50.02 1.1975 ;
      RECT 49.77 0.3075 49.835 0.3725 ;
      RECT 49.77 1.1325 49.835 1.1975 ;
      RECT 49.1825 0.3075 49.2475 0.3725 ;
      RECT 49.1825 1.1325 49.2475 1.1975 ;
      RECT 48.9975 0.3075 49.0625 0.3725 ;
      RECT 48.9975 0.6925 49.0625 0.7575 ;
      RECT 48.9975 1.1325 49.0625 1.1975 ;
      RECT 48.525 0.3075 48.59 0.3725 ;
      RECT 48.525 1.1325 48.59 1.1975 ;
      RECT 48.34 0.3075 48.405 0.3725 ;
      RECT 48.34 0.6825 48.405 0.7475 ;
      RECT 48.34 1.1325 48.405 1.1975 ;
      RECT 48.065 0.6575 48.13 0.7225 ;
      RECT 47.695 0.3075 47.76 0.3725 ;
      RECT 47.54 0.875 47.605 0.94 ;
      RECT 47.2325 0.3075 47.2975 0.3725 ;
      RECT 47.2325 1.1325 47.2975 1.1975 ;
      RECT 47.0475 0.3075 47.1125 0.3725 ;
      RECT 47.0475 1.1325 47.1125 1.1975 ;
      RECT 46.8625 0.3075 46.9275 0.3725 ;
      RECT 46.8625 1.1325 46.9275 1.1975 ;
      RECT 46.275 0.3075 46.34 0.3725 ;
      RECT 46.275 1.1325 46.34 1.1975 ;
      RECT 46.09 0.3075 46.155 0.3725 ;
      RECT 46.09 0.6925 46.155 0.7575 ;
      RECT 46.09 1.1325 46.155 1.1975 ;
      RECT 45.6175 0.3075 45.6825 0.3725 ;
      RECT 45.6175 1.1325 45.6825 1.1975 ;
      RECT 45.4325 0.3075 45.4975 0.3725 ;
      RECT 45.4325 0.6825 45.4975 0.7475 ;
      RECT 45.4325 1.1325 45.4975 1.1975 ;
      RECT 45.1575 0.6575 45.2225 0.7225 ;
      RECT 44.7875 0.3075 44.8525 0.3725 ;
      RECT 44.6325 0.875 44.6975 0.94 ;
      RECT 44.325 0.3075 44.39 0.3725 ;
      RECT 44.325 1.1325 44.39 1.1975 ;
      RECT 44.14 0.3075 44.205 0.3725 ;
      RECT 44.14 1.1325 44.205 1.1975 ;
      RECT 43.955 0.3075 44.02 0.3725 ;
      RECT 43.955 1.1325 44.02 1.1975 ;
      RECT 43.3675 0.3075 43.4325 0.3725 ;
      RECT 43.3675 1.1325 43.4325 1.1975 ;
      RECT 43.1825 0.3075 43.2475 0.3725 ;
      RECT 43.1825 0.6925 43.2475 0.7575 ;
      RECT 43.1825 1.1325 43.2475 1.1975 ;
      RECT 42.71 0.3075 42.775 0.3725 ;
      RECT 42.71 1.1325 42.775 1.1975 ;
      RECT 42.525 0.3075 42.59 0.3725 ;
      RECT 42.525 0.6825 42.59 0.7475 ;
      RECT 42.525 1.1325 42.59 1.1975 ;
      RECT 42.25 0.6575 42.315 0.7225 ;
      RECT 41.88 0.3075 41.945 0.3725 ;
      RECT 41.725 0.875 41.79 0.94 ;
      RECT 41.4175 0.3075 41.4825 0.3725 ;
      RECT 41.4175 1.1325 41.4825 1.1975 ;
      RECT 41.2325 0.3075 41.2975 0.3725 ;
      RECT 41.2325 1.1325 41.2975 1.1975 ;
      RECT 41.0475 0.3075 41.1125 0.3725 ;
      RECT 41.0475 1.1325 41.1125 1.1975 ;
      RECT 40.46 0.3075 40.525 0.3725 ;
      RECT 40.46 1.1325 40.525 1.1975 ;
      RECT 40.275 0.3075 40.34 0.3725 ;
      RECT 40.275 0.6925 40.34 0.7575 ;
      RECT 40.275 1.1325 40.34 1.1975 ;
      RECT 39.8025 0.3075 39.8675 0.3725 ;
      RECT 39.8025 1.1325 39.8675 1.1975 ;
      RECT 39.6175 0.3075 39.6825 0.3725 ;
      RECT 39.6175 0.6825 39.6825 0.7475 ;
      RECT 39.6175 1.1325 39.6825 1.1975 ;
      RECT 39.3425 0.6575 39.4075 0.7225 ;
      RECT 38.9725 0.3075 39.0375 0.3725 ;
      RECT 38.8175 0.875 38.8825 0.94 ;
      RECT 38.51 0.3075 38.575 0.3725 ;
      RECT 38.51 1.1325 38.575 1.1975 ;
      RECT 38.325 0.3075 38.39 0.3725 ;
      RECT 38.325 1.1325 38.39 1.1975 ;
      RECT 38.14 0.3075 38.205 0.3725 ;
      RECT 38.14 1.1325 38.205 1.1975 ;
      RECT 37.5525 0.3075 37.6175 0.3725 ;
      RECT 37.5525 1.1325 37.6175 1.1975 ;
      RECT 37.3675 0.3075 37.4325 0.3725 ;
      RECT 37.3675 0.6925 37.4325 0.7575 ;
      RECT 37.3675 1.1325 37.4325 1.1975 ;
      RECT 36.895 0.3075 36.96 0.3725 ;
      RECT 36.895 1.1325 36.96 1.1975 ;
      RECT 36.71 0.3075 36.775 0.3725 ;
      RECT 36.71 0.6825 36.775 0.7475 ;
      RECT 36.71 1.1325 36.775 1.1975 ;
      RECT 36.435 0.6575 36.5 0.7225 ;
      RECT 36.065 0.3075 36.13 0.3725 ;
      RECT 35.91 0.875 35.975 0.94 ;
      RECT 35.6025 0.3075 35.6675 0.3725 ;
      RECT 35.6025 1.1325 35.6675 1.1975 ;
      RECT 35.4175 0.3075 35.4825 0.3725 ;
      RECT 35.4175 1.1325 35.4825 1.1975 ;
      RECT 35.2325 0.3075 35.2975 0.3725 ;
      RECT 35.2325 1.1325 35.2975 1.1975 ;
      RECT 34.645 0.3075 34.71 0.3725 ;
      RECT 34.645 1.1325 34.71 1.1975 ;
      RECT 34.46 0.3075 34.525 0.3725 ;
      RECT 34.46 0.6925 34.525 0.7575 ;
      RECT 34.46 1.1325 34.525 1.1975 ;
      RECT 33.9875 0.3075 34.0525 0.3725 ;
      RECT 33.9875 1.1325 34.0525 1.1975 ;
      RECT 33.8025 0.3075 33.8675 0.3725 ;
      RECT 33.8025 0.6825 33.8675 0.7475 ;
      RECT 33.8025 1.1325 33.8675 1.1975 ;
      RECT 33.5275 0.6575 33.5925 0.7225 ;
      RECT 33.1575 0.3075 33.2225 0.3725 ;
      RECT 33.0025 0.875 33.0675 0.94 ;
      RECT 32.695 0.3075 32.76 0.3725 ;
      RECT 32.695 1.1325 32.76 1.1975 ;
      RECT 32.51 0.3075 32.575 0.3725 ;
      RECT 32.51 1.1325 32.575 1.1975 ;
      RECT 32.325 0.3075 32.39 0.3725 ;
      RECT 32.325 1.1325 32.39 1.1975 ;
      RECT 31.7375 0.3075 31.8025 0.3725 ;
      RECT 31.7375 1.1325 31.8025 1.1975 ;
      RECT 31.5525 0.3075 31.6175 0.3725 ;
      RECT 31.5525 0.6925 31.6175 0.7575 ;
      RECT 31.5525 1.1325 31.6175 1.1975 ;
      RECT 31.08 0.3075 31.145 0.3725 ;
      RECT 31.08 1.1325 31.145 1.1975 ;
      RECT 30.895 0.3075 30.96 0.3725 ;
      RECT 30.895 0.6825 30.96 0.7475 ;
      RECT 30.895 1.1325 30.96 1.1975 ;
      RECT 30.62 0.6575 30.685 0.7225 ;
      RECT 30.25 0.3075 30.315 0.3725 ;
      RECT 30.095 0.875 30.16 0.94 ;
      RECT 29.7875 0.3075 29.8525 0.3725 ;
      RECT 29.7875 1.1325 29.8525 1.1975 ;
      RECT 29.6025 0.3075 29.6675 0.3725 ;
      RECT 29.6025 1.1325 29.6675 1.1975 ;
      RECT 29.4175 0.3075 29.4825 0.3725 ;
      RECT 29.4175 1.1325 29.4825 1.1975 ;
      RECT 28.83 0.3075 28.895 0.3725 ;
      RECT 28.83 1.1325 28.895 1.1975 ;
      RECT 28.645 0.3075 28.71 0.3725 ;
      RECT 28.645 0.6925 28.71 0.7575 ;
      RECT 28.645 1.1325 28.71 1.1975 ;
      RECT 28.1725 0.3075 28.2375 0.3725 ;
      RECT 28.1725 1.1325 28.2375 1.1975 ;
      RECT 27.9875 0.3075 28.0525 0.3725 ;
      RECT 27.9875 0.6825 28.0525 0.7475 ;
      RECT 27.9875 1.1325 28.0525 1.1975 ;
      RECT 27.7125 0.6575 27.7775 0.7225 ;
      RECT 27.3425 0.3075 27.4075 0.3725 ;
      RECT 27.1875 0.875 27.2525 0.94 ;
      RECT 26.88 0.3075 26.945 0.3725 ;
      RECT 26.88 1.1325 26.945 1.1975 ;
      RECT 26.695 0.3075 26.76 0.3725 ;
      RECT 26.695 1.1325 26.76 1.1975 ;
      RECT 26.51 0.3075 26.575 0.3725 ;
      RECT 26.51 1.1325 26.575 1.1975 ;
      RECT 25.9225 0.3075 25.9875 0.3725 ;
      RECT 25.9225 1.1325 25.9875 1.1975 ;
      RECT 25.7375 0.3075 25.8025 0.3725 ;
      RECT 25.7375 0.6925 25.8025 0.7575 ;
      RECT 25.7375 1.1325 25.8025 1.1975 ;
      RECT 25.265 0.3075 25.33 0.3725 ;
      RECT 25.265 1.1325 25.33 1.1975 ;
      RECT 25.08 0.3075 25.145 0.3725 ;
      RECT 25.08 0.6825 25.145 0.7475 ;
      RECT 25.08 1.1325 25.145 1.1975 ;
      RECT 24.805 0.6575 24.87 0.7225 ;
      RECT 24.435 0.3075 24.5 0.3725 ;
      RECT 24.28 0.875 24.345 0.94 ;
      RECT 23.9725 0.3075 24.0375 0.3725 ;
      RECT 23.9725 1.1325 24.0375 1.1975 ;
      RECT 23.7875 0.3075 23.8525 0.3725 ;
      RECT 23.7875 1.1325 23.8525 1.1975 ;
      RECT 23.6025 0.3075 23.6675 0.3725 ;
      RECT 23.6025 1.1325 23.6675 1.1975 ;
      RECT 23.015 0.3075 23.08 0.3725 ;
      RECT 23.015 1.1325 23.08 1.1975 ;
      RECT 22.83 0.3075 22.895 0.3725 ;
      RECT 22.83 0.6925 22.895 0.7575 ;
      RECT 22.83 1.1325 22.895 1.1975 ;
      RECT 22.3575 0.3075 22.4225 0.3725 ;
      RECT 22.3575 1.1325 22.4225 1.1975 ;
      RECT 22.1725 0.3075 22.2375 0.3725 ;
      RECT 22.1725 0.6825 22.2375 0.7475 ;
      RECT 22.1725 1.1325 22.2375 1.1975 ;
      RECT 21.8975 0.6575 21.9625 0.7225 ;
      RECT 21.5275 0.3075 21.5925 0.3725 ;
      RECT 21.3725 0.875 21.4375 0.94 ;
      RECT 21.065 0.3075 21.13 0.3725 ;
      RECT 21.065 1.1325 21.13 1.1975 ;
      RECT 20.88 0.3075 20.945 0.3725 ;
      RECT 20.88 1.1325 20.945 1.1975 ;
      RECT 20.695 0.3075 20.76 0.3725 ;
      RECT 20.695 1.1325 20.76 1.1975 ;
      RECT 20.1075 0.3075 20.1725 0.3725 ;
      RECT 20.1075 1.1325 20.1725 1.1975 ;
      RECT 19.9225 0.3075 19.9875 0.3725 ;
      RECT 19.9225 0.6925 19.9875 0.7575 ;
      RECT 19.9225 1.1325 19.9875 1.1975 ;
      RECT 19.45 0.3075 19.515 0.3725 ;
      RECT 19.45 1.1325 19.515 1.1975 ;
      RECT 19.265 0.3075 19.33 0.3725 ;
      RECT 19.265 0.6825 19.33 0.7475 ;
      RECT 19.265 1.1325 19.33 1.1975 ;
      RECT 18.99 0.6575 19.055 0.7225 ;
      RECT 18.62 0.3075 18.685 0.3725 ;
      RECT 18.465 0.875 18.53 0.94 ;
      RECT 18.1575 0.3075 18.2225 0.3725 ;
      RECT 18.1575 1.1325 18.2225 1.1975 ;
      RECT 17.9725 0.3075 18.0375 0.3725 ;
      RECT 17.9725 1.1325 18.0375 1.1975 ;
      RECT 17.7875 0.3075 17.8525 0.3725 ;
      RECT 17.7875 1.1325 17.8525 1.1975 ;
      RECT 17.2 0.3075 17.265 0.3725 ;
      RECT 17.2 1.1325 17.265 1.1975 ;
      RECT 17.015 0.3075 17.08 0.3725 ;
      RECT 17.015 0.6925 17.08 0.7575 ;
      RECT 17.015 1.1325 17.08 1.1975 ;
      RECT 16.5425 0.3075 16.6075 0.3725 ;
      RECT 16.5425 1.1325 16.6075 1.1975 ;
      RECT 16.3575 0.3075 16.4225 0.3725 ;
      RECT 16.3575 0.6825 16.4225 0.7475 ;
      RECT 16.3575 1.1325 16.4225 1.1975 ;
      RECT 16.0825 0.6575 16.1475 0.7225 ;
      RECT 15.7125 0.3075 15.7775 0.3725 ;
      RECT 15.5575 0.875 15.6225 0.94 ;
      RECT 15.25 0.3075 15.315 0.3725 ;
      RECT 15.25 1.1325 15.315 1.1975 ;
      RECT 15.065 0.3075 15.13 0.3725 ;
      RECT 15.065 1.1325 15.13 1.1975 ;
      RECT 14.88 0.3075 14.945 0.3725 ;
      RECT 14.88 1.1325 14.945 1.1975 ;
      RECT 14.2925 0.3075 14.3575 0.3725 ;
      RECT 14.2925 1.1325 14.3575 1.1975 ;
      RECT 14.1075 0.3075 14.1725 0.3725 ;
      RECT 14.1075 0.6925 14.1725 0.7575 ;
      RECT 14.1075 1.1325 14.1725 1.1975 ;
      RECT 13.635 0.3075 13.7 0.3725 ;
      RECT 13.635 1.1325 13.7 1.1975 ;
      RECT 13.45 0.3075 13.515 0.3725 ;
      RECT 13.45 0.6825 13.515 0.7475 ;
      RECT 13.45 1.1325 13.515 1.1975 ;
      RECT 13.175 0.6575 13.24 0.7225 ;
      RECT 12.805 0.3075 12.87 0.3725 ;
      RECT 12.65 0.875 12.715 0.94 ;
      RECT 12.3425 0.3075 12.4075 0.3725 ;
      RECT 12.3425 1.1325 12.4075 1.1975 ;
      RECT 12.1575 0.3075 12.2225 0.3725 ;
      RECT 12.1575 1.1325 12.2225 1.1975 ;
      RECT 11.9725 0.3075 12.0375 0.3725 ;
      RECT 11.9725 1.1325 12.0375 1.1975 ;
      RECT 11.385 0.3075 11.45 0.3725 ;
      RECT 11.385 1.1325 11.45 1.1975 ;
      RECT 11.2 0.3075 11.265 0.3725 ;
      RECT 11.2 0.6925 11.265 0.7575 ;
      RECT 11.2 1.1325 11.265 1.1975 ;
      RECT 10.7275 0.3075 10.7925 0.3725 ;
      RECT 10.7275 1.1325 10.7925 1.1975 ;
      RECT 10.5425 0.3075 10.6075 0.3725 ;
      RECT 10.5425 0.6825 10.6075 0.7475 ;
      RECT 10.5425 1.1325 10.6075 1.1975 ;
      RECT 10.2675 0.6575 10.3325 0.7225 ;
      RECT 9.8975 0.3075 9.9625 0.3725 ;
      RECT 9.7425 0.875 9.8075 0.94 ;
      RECT 9.435 0.3075 9.5 0.3725 ;
      RECT 9.435 1.1325 9.5 1.1975 ;
      RECT 9.25 0.3075 9.315 0.3725 ;
      RECT 9.25 1.1325 9.315 1.1975 ;
      RECT 9.065 0.3075 9.13 0.3725 ;
      RECT 9.065 1.1325 9.13 1.1975 ;
      RECT 8.4775 0.3075 8.5425 0.3725 ;
      RECT 8.4775 1.1325 8.5425 1.1975 ;
      RECT 8.2925 0.3075 8.3575 0.3725 ;
      RECT 8.2925 0.6925 8.3575 0.7575 ;
      RECT 8.2925 1.1325 8.3575 1.1975 ;
      RECT 7.82 0.3075 7.885 0.3725 ;
      RECT 7.82 1.1325 7.885 1.1975 ;
      RECT 7.635 0.3075 7.7 0.3725 ;
      RECT 7.635 0.6825 7.7 0.7475 ;
      RECT 7.635 1.1325 7.7 1.1975 ;
      RECT 7.36 0.6575 7.425 0.7225 ;
      RECT 6.99 0.3075 7.055 0.3725 ;
      RECT 6.835 0.875 6.9 0.94 ;
      RECT 6.5275 0.3075 6.5925 0.3725 ;
      RECT 6.5275 1.1325 6.5925 1.1975 ;
      RECT 6.3425 0.3075 6.4075 0.3725 ;
      RECT 6.3425 1.1325 6.4075 1.1975 ;
      RECT 6.1575 0.3075 6.2225 0.3725 ;
      RECT 6.1575 1.1325 6.2225 1.1975 ;
      RECT 5.57 0.3075 5.635 0.3725 ;
      RECT 5.57 1.1325 5.635 1.1975 ;
      RECT 5.385 0.3075 5.45 0.3725 ;
      RECT 5.385 0.6925 5.45 0.7575 ;
      RECT 5.385 1.1325 5.45 1.1975 ;
      RECT 4.9125 0.3075 4.9775 0.3725 ;
      RECT 4.9125 1.1325 4.9775 1.1975 ;
      RECT 4.7275 0.3075 4.7925 0.3725 ;
      RECT 4.7275 0.6825 4.7925 0.7475 ;
      RECT 4.7275 1.1325 4.7925 1.1975 ;
      RECT 4.4525 0.6575 4.5175 0.7225 ;
      RECT 4.0825 0.3075 4.1475 0.3725 ;
      RECT 3.9275 0.875 3.9925 0.94 ;
      RECT 3.62 0.3075 3.685 0.3725 ;
      RECT 3.62 1.1325 3.685 1.1975 ;
      RECT 3.435 0.3075 3.5 0.3725 ;
      RECT 3.435 1.1325 3.5 1.1975 ;
      RECT 3.25 0.3075 3.315 0.3725 ;
      RECT 3.25 1.1325 3.315 1.1975 ;
      RECT 2.6625 0.3075 2.7275 0.3725 ;
      RECT 2.6625 1.1325 2.7275 1.1975 ;
      RECT 2.4775 0.3075 2.5425 0.3725 ;
      RECT 2.4775 0.6925 2.5425 0.7575 ;
      RECT 2.4775 1.1325 2.5425 1.1975 ;
      RECT 2.005 0.3075 2.07 0.3725 ;
      RECT 2.005 1.1325 2.07 1.1975 ;
      RECT 1.82 0.3075 1.885 0.3725 ;
      RECT 1.82 0.6825 1.885 0.7475 ;
      RECT 1.82 1.1325 1.885 1.1975 ;
      RECT 1.545 0.6575 1.61 0.7225 ;
      RECT 1.175 0.3075 1.24 0.3725 ;
      RECT 1.02 0.875 1.085 0.94 ;
      RECT 0.7125 0.3075 0.7775 0.3725 ;
      RECT 0.7125 1.1325 0.7775 1.1975 ;
      RECT 0.5275 0.3075 0.5925 0.3725 ;
      RECT 0.5275 1.1325 0.5925 1.1975 ;
      RECT 0.3425 0.3075 0.4075 0.3725 ;
      RECT 0.3425 1.1325 0.4075 1.1975 ;
    LAYER via2 ;
      RECT 93.8575 0.785 93.9275 0.855 ;
      RECT 91.8275 0.785 91.8975 0.855 ;
      RECT 91.4925 1.13 91.5625 1.2 ;
      RECT 90.835 0.305 90.905 0.375 ;
      RECT 89.885 1.13 89.955 1.2 ;
      RECT 89.2275 0.305 89.2975 0.375 ;
      RECT 86.9775 1.13 87.0475 1.2 ;
      RECT 86.32 0.305 86.39 0.375 ;
      RECT 84.07 1.13 84.14 1.2 ;
      RECT 83.4125 0.305 83.4825 0.375 ;
      RECT 81.1625 1.13 81.2325 1.2 ;
      RECT 80.505 0.305 80.575 0.375 ;
      RECT 78.255 1.13 78.325 1.2 ;
      RECT 77.5975 0.305 77.6675 0.375 ;
      RECT 75.3475 1.13 75.4175 1.2 ;
      RECT 74.69 0.305 74.76 0.375 ;
      RECT 72.44 1.13 72.51 1.2 ;
      RECT 71.7825 0.305 71.8525 0.375 ;
      RECT 69.5325 1.13 69.6025 1.2 ;
      RECT 68.875 0.305 68.945 0.375 ;
      RECT 66.625 1.13 66.695 1.2 ;
      RECT 65.9675 0.305 66.0375 0.375 ;
      RECT 63.7175 1.13 63.7875 1.2 ;
      RECT 63.06 0.305 63.13 0.375 ;
      RECT 60.81 1.13 60.88 1.2 ;
      RECT 60.1525 0.305 60.2225 0.375 ;
      RECT 57.9025 1.13 57.9725 1.2 ;
      RECT 57.245 0.305 57.315 0.375 ;
      RECT 54.995 1.13 55.065 1.2 ;
      RECT 54.3375 0.305 54.4075 0.375 ;
      RECT 52.0875 1.13 52.1575 1.2 ;
      RECT 51.43 0.305 51.5 0.375 ;
      RECT 49.18 1.13 49.25 1.2 ;
      RECT 48.5225 0.305 48.5925 0.375 ;
      RECT 46.2725 1.13 46.3425 1.2 ;
      RECT 45.615 0.305 45.685 0.375 ;
      RECT 43.365 1.13 43.435 1.2 ;
      RECT 42.7075 0.305 42.7775 0.375 ;
      RECT 40.4575 1.13 40.5275 1.2 ;
      RECT 39.8 0.305 39.87 0.375 ;
      RECT 37.55 1.13 37.62 1.2 ;
      RECT 36.8925 0.305 36.9625 0.375 ;
      RECT 34.6425 1.13 34.7125 1.2 ;
      RECT 33.985 0.305 34.055 0.375 ;
      RECT 31.735 1.13 31.805 1.2 ;
      RECT 31.0775 0.305 31.1475 0.375 ;
      RECT 28.8275 1.13 28.8975 1.2 ;
      RECT 28.17 0.305 28.24 0.375 ;
      RECT 25.92 1.13 25.99 1.2 ;
      RECT 25.2625 0.305 25.3325 0.375 ;
      RECT 23.0125 1.13 23.0825 1.2 ;
      RECT 22.355 0.305 22.425 0.375 ;
      RECT 20.105 1.13 20.175 1.2 ;
      RECT 19.4475 0.305 19.5175 0.375 ;
      RECT 17.1975 1.13 17.2675 1.2 ;
      RECT 16.54 0.305 16.61 0.375 ;
      RECT 14.29 1.13 14.36 1.2 ;
      RECT 13.6325 0.305 13.7025 0.375 ;
      RECT 11.3825 1.13 11.4525 1.2 ;
      RECT 10.725 0.305 10.795 0.375 ;
      RECT 8.475 1.13 8.545 1.2 ;
      RECT 7.8175 0.305 7.8875 0.375 ;
      RECT 5.5675 1.13 5.6375 1.2 ;
      RECT 4.91 0.305 4.98 0.375 ;
      RECT 2.66 1.13 2.73 1.2 ;
      RECT 2.0025 0.305 2.0725 0.375 ;
    LAYER via3 ;
      RECT 93.8575 0.785 93.9275 0.855 ;
      RECT 91.8275 0.785 91.8975 0.855 ;
      RECT 91.4925 1.13 91.5625 1.2 ;
      RECT 90.835 0.305 90.905 0.375 ;
      RECT 89.885 1.13 89.955 1.2 ;
      RECT 89.2275 0.305 89.2975 0.375 ;
      RECT 86.9775 1.13 87.0475 1.2 ;
      RECT 86.32 0.305 86.39 0.375 ;
      RECT 84.07 1.13 84.14 1.2 ;
      RECT 83.4125 0.305 83.4825 0.375 ;
      RECT 81.1625 1.13 81.2325 1.2 ;
      RECT 80.505 0.305 80.575 0.375 ;
      RECT 78.255 1.13 78.325 1.2 ;
      RECT 77.5975 0.305 77.6675 0.375 ;
      RECT 75.3475 1.13 75.4175 1.2 ;
      RECT 74.69 0.305 74.76 0.375 ;
      RECT 72.44 1.13 72.51 1.2 ;
      RECT 71.7825 0.305 71.8525 0.375 ;
      RECT 69.5325 1.13 69.6025 1.2 ;
      RECT 68.875 0.305 68.945 0.375 ;
      RECT 66.625 1.13 66.695 1.2 ;
      RECT 65.9675 0.305 66.0375 0.375 ;
      RECT 63.7175 1.13 63.7875 1.2 ;
      RECT 63.06 0.305 63.13 0.375 ;
      RECT 60.81 1.13 60.88 1.2 ;
      RECT 60.1525 0.305 60.2225 0.375 ;
      RECT 57.9025 1.13 57.9725 1.2 ;
      RECT 57.245 0.305 57.315 0.375 ;
      RECT 54.995 1.13 55.065 1.2 ;
      RECT 54.3375 0.305 54.4075 0.375 ;
      RECT 52.0875 1.13 52.1575 1.2 ;
      RECT 51.43 0.305 51.5 0.375 ;
      RECT 49.18 1.13 49.25 1.2 ;
      RECT 48.5225 0.305 48.5925 0.375 ;
      RECT 46.2725 1.13 46.3425 1.2 ;
      RECT 45.615 0.305 45.685 0.375 ;
      RECT 43.365 1.13 43.435 1.2 ;
      RECT 42.7075 0.305 42.7775 0.375 ;
      RECT 40.4575 1.13 40.5275 1.2 ;
      RECT 39.8 0.305 39.87 0.375 ;
      RECT 37.55 1.13 37.62 1.2 ;
      RECT 36.8925 0.305 36.9625 0.375 ;
      RECT 34.6425 1.13 34.7125 1.2 ;
      RECT 33.985 0.305 34.055 0.375 ;
      RECT 31.735 1.13 31.805 1.2 ;
      RECT 31.0775 0.305 31.1475 0.375 ;
      RECT 28.8275 1.13 28.8975 1.2 ;
      RECT 28.17 0.305 28.24 0.375 ;
      RECT 25.92 1.13 25.99 1.2 ;
      RECT 25.2625 0.305 25.3325 0.375 ;
      RECT 23.0125 1.13 23.0825 1.2 ;
      RECT 22.355 0.305 22.425 0.375 ;
      RECT 20.105 1.13 20.175 1.2 ;
      RECT 19.4475 0.305 19.5175 0.375 ;
      RECT 17.1975 1.13 17.2675 1.2 ;
      RECT 16.54 0.305 16.61 0.375 ;
      RECT 14.29 1.13 14.36 1.2 ;
      RECT 13.6325 0.305 13.7025 0.375 ;
      RECT 11.3825 1.13 11.4525 1.2 ;
      RECT 10.725 0.305 10.795 0.375 ;
      RECT 8.475 1.13 8.545 1.2 ;
      RECT 7.8175 0.305 7.8875 0.375 ;
      RECT 5.5675 1.13 5.6375 1.2 ;
      RECT 4.91 0.305 4.98 0.375 ;
      RECT 2.66 1.13 2.73 1.2 ;
      RECT 2.0025 0.305 2.0725 0.375 ;
  END
END regfile

END LIBRARY
