/home/soumilg2/Documents/ece425_work/mp_pnr/provided/regfile.lef