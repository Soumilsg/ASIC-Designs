VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER contactResistance REAL ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.0025 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER contact
  TYPE CUT ;
  SPACING 0.075 ;
  PROPERTY contactResistance 10.5 ;
END contact

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.065 ;
  SPACING 0.065 ;
  SPACING 0.065 SAMENET ;
  RESISTANCE RPERSQ 0.38 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.065 ;
  PROPERTY contactResistance 5.69 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.075 ;
  SPACING 0.07 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
  PROPERTY contactResistance 11.39 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.07 ;
  SPACING 0.07 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
  PROPERTY contactResistance 16.73 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 21.44 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal5

LAYER via5
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 24.08 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal6

LAYER via6
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 11.39 ;
END via6

LAYER metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.855 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.44 ;
  SPACING 0.44 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal7

LAYER via7
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  PROPERTY contactResistance 5.69 ;
END via7

LAYER metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.855 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.44 ;
  SPACING 0.44 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal8

LAYER via8
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  PROPERTY contactResistance 16.73 ;
END via8

LAYER metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.71 1.71 ;
  WIDTH 0.8 ;
  SPACING 0.8 ;
  SPACING 0.8 SAMENET ;
  RESISTANCE RPERSQ 0.21 ;
END metal9

LAYER via9
  TYPE CUT ;
  SPACING 0.88 ;
  WIDTH 0.8 ;
  PROPERTY contactResistance 21.44 ;
END via9

LAYER metal10
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.71 1.71 ;
  WIDTH 0.4 ;
  SPACING 0.8 ;
  SPACING 0.8 SAMENET ;
  RESISTANCE RPERSQ 0.21 ;
END metal10

VIARULE M2_M1 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M2_M1

VIARULE M3_M2 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M3_M2

VIARULE M4_M3 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M4_M3

VIARULE M5_M4 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M5_M4

VIARULE M6_M5 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M6_M5

VIARULE M7_M6 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M7_M6

VIARULE M8_M7 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 0.8 ;
END M8_M7

VIARULE M9_M8 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 0.8 ;
END M9_M8

VIARULE M10_M9 GENERATE
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.6 BY 1.6 ;
END M10_M9

VIARULE M1_POLY GENERATE
  LAYER poly ;
    ENCLOSURE 0 0 ;
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER contact ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M1_POLY

VIA M2_M1_via DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_via

VIA M3_M2_via DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_via

VIA M4_M3_via DEFAULT
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_via

VIA M5_M4_via DEFAULT
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M5_M4_via

VIA M6_M5_via DEFAULT
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M6_M5_via

VIA M7_M6_via DEFAULT
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M7_M6_via

VIA M8_M7_via DEFAULT
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M8_M7_via

VIA M9_M8_via DEFAULT
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M9_M8_via

VIA M10_M9_via DEFAULT
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal10 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M10_M9_via

VIA M2_M1_viaB DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.0675 -0.035 0.0675 0.035 ;
END M2_M1_viaB

VIA M2_M1_viaC DEFAULT
  LAYER metal1 ;
    RECT -0.0325 -0.0675 0.0325 0.0675 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_viaC

VIA M3_M2_viaB DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END M3_M2_viaB

VIA M3_M2_viaC DEFAULT
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_viaC

VIA M4_M3_viaB DEFAULT
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_viaB

SITE CoreSite
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.005 BY 1.005 ;
END CoreSite

MACRO and2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN and2 0 0.1 ;
  SIZE 0.75 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1975 0.4625 0.2625 0.5975 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.275 0.6625 0.41 0.7275 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.625 0.265 0.69 1.2825 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 0.745 1.55 ;
        RECT 0.435 1.0425 0.5 1.55 ;
        RECT 0.06 1.04 0.125 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.75 0.2 ;
        RECT 0.435 0 0.5 0.415 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.2475 0.825 0.3125 1.2825 ;
      RECT 0.48 0.79 0.545 0.925 ;
      RECT 0.06 0.825 0.545 0.89 ;
      RECT 0.06 0.265 0.125 0.89 ;
  END
END and2

MACRO aoi21
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN aoi21 0 0.1 ;
  SIZE 0.75 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.09 0.8175 0.155 0.9525 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.29 0.8175 0.355 0.9525 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.48 0.8175 0.545 0.9525 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.625 0.265 0.69 1.2825 ;
        RECT 0.06 0.5575 0.69 0.6225 ;
        RECT 0.06 0.265 0.125 0.6225 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 0.755 1.55 ;
        RECT 0.2475 1.04 0.3125 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.75 0.2 ;
        RECT 0.435 0 0.5 0.415 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.435 1.0525 0.5 1.2725 ;
      RECT 0.06 1.0525 0.125 1.2725 ;
    LAYER metal2 ;
      RECT 0.0575 1.2925 0.5025 1.3625 ;
      RECT 0.4325 1.0975 0.5025 1.3625 ;
      RECT 0.0575 1.0975 0.1275 1.3625 ;
    LAYER via1 ;
      RECT 0.435 1.1325 0.5 1.1975 ;
      RECT 0.06 1.1325 0.125 1.1975 ;
  END
END aoi21

MACRO buf
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN buf 0 0.1 ;
  SIZE 0.56 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2025 0.7075 0.2675 0.8425 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.435 0.265 0.5 1.285 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 0.56 1.55 ;
        RECT 0.245 1.045 0.31 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.56 0.2 ;
        RECT 0.245 0 0.31 0.4225 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.06 0.265 0.125 1.285 ;
      RECT 0.2925 0.505 0.3575 0.64 ;
      RECT 0.06 0.54 0.3575 0.605 ;
  END
END buf

MACRO dff
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN dff 0 0.1 ;
  SIZE 3.7 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.7875 0.18 0.8525 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.575 0.265 3.64 1.285 ;
        RECT 3.15 0.53 3.64 0.595 ;
    END
  END Q
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 3.7 1.55 ;
        RECT 3.39 1.045 3.455 1.55 ;
        RECT 3.205 1.045 3.27 1.55 ;
        RECT 1.91 1.045 1.975 1.55 ;
        RECT 1.725 1.045 1.79 1.55 ;
        RECT 0.43 1.045 0.495 1.55 ;
        RECT 0.06 1.045 0.125 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 3.7 0.2 ;
        RECT 3.39 0 3.455 0.4225 ;
        RECT 3.205 0 3.27 0.4225 ;
        RECT 1.91 0 1.975 0.4225 ;
        RECT 1.725 0 1.79 0.4225 ;
        RECT 0.43 0 0.495 0.4225 ;
        RECT 0.06 0 0.125 0.4225 ;
    END
  END vss!
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.7975 0.2725 0.8675 1.235 ;
      LAYER metal1 ;
        RECT 0.8 0.265 0.865 0.415 ;
        RECT 0.8 1.045 0.865 1.285 ;
      LAYER via1 ;
        RECT 0.8 1.135 0.865 1.2 ;
        RECT 0.8 0.3075 0.865 0.3725 ;
    END
  END D
  OBS
    LAYER metal1 ;
      RECT 0.245 0.265 0.31 1.285 ;
      RECT 0.245 0.91 2.4725 0.975 ;
      RECT 2.37 0.7375 2.435 0.975 ;
      RECT 2.37 0.7375 2.8075 0.8025 ;
      RECT 2.7425 0.5275 2.8075 0.8025 ;
      RECT 0.245 0.6275 0.5375 0.6925 ;
      RECT 2.7075 0.5275 2.8425 0.5925 ;
      RECT 0.245 0.4925 0.9925 0.5575 ;
      RECT 2.095 0.4975 2.16 0.6325 ;
      RECT 1.67 0.5325 2.16 0.5975 ;
      RECT 0.58 0.775 1.3275 0.84 ;
      RECT 1.2625 0.5275 1.3275 0.84 ;
      RECT 1.2275 0.5275 1.3625 0.5925 ;
      RECT 3.375 0.7875 3.51 0.8525 ;
      RECT 3.02 0.265 3.085 1.285 ;
      RECT 2.835 0.265 2.9 0.415 ;
      RECT 2.835 1.045 2.9 1.285 ;
      RECT 2.65 0.265 2.715 0.415 ;
      RECT 2.65 1.045 2.715 1.285 ;
      RECT 2.465 0.265 2.53 0.415 ;
      RECT 2.465 1.045 2.53 1.285 ;
      RECT 2.28 0.265 2.345 0.415 ;
      RECT 2.28 1.045 2.345 1.285 ;
      RECT 2.095 0.265 2.16 0.415 ;
      RECT 2.095 1.045 2.16 1.285 ;
      RECT 1.93 0.7025 1.995 0.8375 ;
      RECT 1.54 0.265 1.605 0.415 ;
      RECT 1.54 1.045 1.605 1.285 ;
      RECT 1.355 0.265 1.42 0.415 ;
      RECT 1.355 1.045 1.42 1.285 ;
      RECT 1.17 0.265 1.235 0.415 ;
      RECT 1.17 1.045 1.235 1.285 ;
      RECT 0.985 0.265 1.05 0.415 ;
      RECT 0.985 1.045 1.05 1.285 ;
      RECT 0.615 0.265 0.68 0.415 ;
      RECT 0.615 1.045 0.68 1.285 ;
    LAYER metal2 ;
      RECT 2.6475 0.125 2.7175 1.235 ;
      RECT 2.4625 0.125 2.5325 1.235 ;
      RECT 3.375 0.785 3.51 0.855 ;
      RECT 3.4075 0.125 3.4775 0.855 ;
      RECT 2.4625 0.125 3.4775 0.195 ;
      RECT 2.8325 0.2725 2.9025 1.235 ;
      RECT 3.0175 0.825 3.0875 0.96 ;
      RECT 2.8325 0.8575 3.0875 0.9275 ;
      RECT 2.2775 0.2725 2.3475 1.235 ;
      RECT 2.0925 0.2725 2.1625 1.235 ;
      RECT 2.0925 0.53 2.3475 0.6 ;
      RECT 1.1675 0.125 1.2375 1.235 ;
      RECT 0.9825 0.125 1.0525 1.235 ;
      RECT 1.9275 0.125 1.9975 0.8375 ;
      RECT 0.9825 0.125 1.9975 0.195 ;
      RECT 1.5375 0.2725 1.6075 1.235 ;
      RECT 1.3525 0.2725 1.4225 1.235 ;
      RECT 1.3525 0.5175 1.6075 0.5875 ;
      RECT 0.6125 0.2725 0.6825 1.285 ;
      RECT 0.58 0.7725 0.715 0.8425 ;
    LAYER via1 ;
      RECT 3.41 0.7875 3.475 0.8525 ;
      RECT 3.02 0.86 3.085 0.925 ;
      RECT 2.835 0.3075 2.9 0.3725 ;
      RECT 2.835 1.135 2.9 1.2 ;
      RECT 2.65 0.3075 2.715 0.3725 ;
      RECT 2.65 1.135 2.715 1.2 ;
      RECT 2.465 0.3075 2.53 0.3725 ;
      RECT 2.465 1.135 2.53 1.2 ;
      RECT 2.28 0.3075 2.345 0.3725 ;
      RECT 2.28 1.135 2.345 1.2 ;
      RECT 2.095 0.3075 2.16 0.3725 ;
      RECT 2.095 0.5325 2.16 0.5975 ;
      RECT 2.095 1.135 2.16 1.2 ;
      RECT 1.93 0.7375 1.995 0.8025 ;
      RECT 1.54 0.3075 1.605 0.3725 ;
      RECT 1.54 1.135 1.605 1.2 ;
      RECT 1.355 0.3075 1.42 0.3725 ;
      RECT 1.355 1.135 1.42 1.2 ;
      RECT 1.17 0.3075 1.235 0.3725 ;
      RECT 1.17 1.135 1.235 1.2 ;
      RECT 0.985 0.3075 1.05 0.3725 ;
      RECT 0.985 1.135 1.05 1.2 ;
      RECT 0.615 0.3075 0.68 0.3725 ;
      RECT 0.615 0.775 0.68 0.84 ;
      RECT 0.615 1.1325 0.68 1.1975 ;
  END
END dff

MACRO inv
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN inv 0 0.1 ;
  SIZE 0.37 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.7875 0.18 0.8525 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.245 0.265 0.31 1.285 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 0.37 1.55 ;
        RECT 0.06 1.045 0.125 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.37 0.2 ;
        RECT 0.06 0 0.125 0.4225 ;
    END
  END vss!
END inv

MACRO latch
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN latch 0 0.1 ;
  SIZE 1.66 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.535 0.265 1.6 1.285 ;
        RECT 1.28 0.5325 1.6 0.5975 ;
        RECT 1.28 0.4975 1.345 0.6325 ;
    END
  END Q
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 1.66 1.55 ;
        RECT 1.345 1.045 1.41 1.55 ;
        RECT 0.59 1.045 0.655 1.55 ;
        RECT 0.245 1.045 0.31 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 1.66 0.2 ;
        RECT 1.345 0 1.41 0.4225 ;
        RECT 0.59 0 0.655 0.4225 ;
        RECT 0.245 0 0.31 0.4225 ;
    END
  END vss!
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.5725 0.7075 0.6425 0.8425 ;
      LAYER metal1 ;
        RECT 0.575 0.7075 0.64 0.8425 ;
      LAYER via1 ;
        RECT 0.575 0.7425 0.64 0.8075 ;
    END
  END D
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.2 0.7075 0.27 0.8425 ;
      LAYER metal1 ;
        RECT 0.2025 0.7075 0.2675 0.8425 ;
      LAYER via1 ;
        RECT 0.2025 0.7425 0.2675 0.8075 ;
    END
  END EN
  OBS
    LAYER metal1 ;
      RECT 0.8725 0.715 0.9375 0.85 ;
      RECT 0.8725 0.75 1.1225 0.815 ;
      RECT 1.0575 0.5125 1.1225 0.815 ;
      RECT 0.435 0.265 0.5 1.285 ;
      RECT 1.0575 0.88 1.1225 1.015 ;
      RECT 0.7375 0.915 1.1225 0.98 ;
      RECT 0.7375 0.55 0.8025 0.98 ;
      RECT 0.8725 0.515 0.9375 0.65 ;
      RECT 0.435 0.5525 0.8025 0.6175 ;
      RECT 0.7375 0.55 0.9375 0.615 ;
      RECT 0.06 0.265 0.125 1.285 ;
      RECT 0.2925 0.505 0.3575 0.64 ;
      RECT 0.06 0.54 0.3575 0.605 ;
      RECT 1.395 0.785 1.46 0.92 ;
      RECT 1.1575 0.2725 1.2225 0.4075 ;
      RECT 1.1575 1.0975 1.2225 1.2325 ;
      RECT 0.965 0.2725 1.03 0.4075 ;
      RECT 0.965 1.0975 1.03 1.2325 ;
      RECT 0.775 0.2725 0.84 0.4075 ;
      RECT 0.775 1.0975 0.84 1.2325 ;
    LAYER metal2 ;
      RECT 0.9625 1.3775 1.4625 1.4475 ;
      RECT 1.3925 0.785 1.4625 1.4475 ;
      RECT 0.9625 0.265 1.0325 1.4475 ;
      RECT 1.155 0.2725 1.225 1.2325 ;
      RECT 0.7725 0.2675 0.8425 1.2325 ;
    LAYER via1 ;
      RECT 1.395 0.82 1.46 0.885 ;
      RECT 1.1575 0.3075 1.2225 0.3725 ;
      RECT 1.1575 1.1325 1.2225 1.1975 ;
      RECT 0.965 0.3075 1.03 0.3725 ;
      RECT 0.965 1.1325 1.03 1.1975 ;
      RECT 0.775 0.3075 0.84 0.3725 ;
      RECT 0.775 1.1325 0.84 1.1975 ;
  END
END latch

MACRO mux2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN mux2 0 0.1 ;
  SIZE 1.32 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.735 0.7425 0.945 0.8125 ;
        RECT 0.875 0.525 0.945 0.8125 ;
        RECT 0.3425 0.525 0.945 0.595 ;
        RECT 0.735 0.71 0.805 0.845 ;
        RECT 0.3075 0.5275 0.4425 0.5975 ;
      LAYER metal1 ;
        RECT 0.7375 0.71 0.8025 0.845 ;
        RECT 0.3075 0.53 0.4425 0.595 ;
      LAYER via1 ;
        RECT 0.3425 0.53 0.4075 0.595 ;
        RECT 0.7375 0.745 0.8025 0.81 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.345 0.95 0.975 1.015 ;
        RECT 0.91 0.575 0.975 1.015 ;
        RECT 0.705 0.575 0.975 0.64 ;
        RECT 0.345 0.71 0.41 1.015 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.195 0.265 1.26 1.285 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 1.32 1.55 ;
        RECT 1.01 1.105 1.075 1.55 ;
        RECT 0.245 1.0825 0.31 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 1.32 0.2 ;
        RECT 1.01 0 1.075 0.505 ;
        RECT 0.245 0 0.31 0.41 ;
    END
  END vss!
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.19 0.74 0.26 0.875 ;
      LAYER metal1 ;
        RECT 0.1925 0.74 0.2575 0.875 ;
      LAYER via1 ;
        RECT 0.1925 0.775 0.2575 0.84 ;
    END
  END S0
  OBS
    LAYER metal1 ;
      RECT 0.06 0.265 0.125 1.285 ;
      RECT 0.0575 0.5475 0.125 0.6825 ;
      RECT 1.0525 0.57 1.1175 0.705 ;
      RECT 0.8175 1.1025 0.8825 1.2375 ;
      RECT 0.6275 0.2675 0.6925 0.4025 ;
      RECT 0.6275 1.13 0.6925 1.265 ;
      RECT 0.4875 0.775 0.6225 0.84 ;
      RECT 0.4375 1.1025 0.5025 1.2375 ;
    LAYER metal2 ;
      RECT 0.625 0.9575 0.695 1.265 ;
      RECT 0.625 0.9575 1.12 1.0275 ;
      RECT 1.05 0.13 1.12 1.0275 ;
      RECT 0.625 0.13 0.695 0.4025 ;
      RECT 0.625 0.13 1.12 0.2 ;
      RECT 0.435 1.375 0.885 1.445 ;
      RECT 0.815 1.1025 0.885 1.445 ;
      RECT 0.435 1.1025 0.505 1.445 ;
      RECT 0.05 0.955 0.555 1.025 ;
      RECT 0.485 0.7725 0.555 1.025 ;
      RECT 0.05 0.5475 0.12 1.025 ;
      RECT 0.485 0.7725 0.6225 0.8425 ;
      RECT 0.05 0.5475 0.125 0.6825 ;
    LAYER via1 ;
      RECT 1.0525 0.605 1.1175 0.67 ;
      RECT 0.8175 1.1375 0.8825 1.2025 ;
      RECT 0.6275 0.3025 0.6925 0.3675 ;
      RECT 0.6275 1.165 0.6925 1.23 ;
      RECT 0.5225 0.775 0.5875 0.84 ;
      RECT 0.4375 1.1375 0.5025 1.2025 ;
      RECT 0.0575 0.5825 0.1225 0.6475 ;
  END
END mux2

MACRO nand2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN nand2 0 0.1 ;
  SIZE 0.56 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1975 0.4975 0.2625 0.6325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.275 0.7525 0.41 0.8175 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.9025 0.56 0.9675 ;
        RECT 0.2475 0.9025 0.3125 1.2825 ;
        RECT 0.06 0.265 0.125 0.9675 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 0.56 1.55 ;
        RECT 0.435 1.0425 0.5 1.55 ;
        RECT 0.06 1.04 0.125 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.56 0.2 ;
        RECT 0.435 0 0.5 0.415 ;
    END
  END vss!
END nand2

MACRO nor2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN nor2 0 0.1 ;
  SIZE 0.56 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.09 0.4975 0.155 0.6325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.38 0.7525 0.515 0.8175 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.245 0.9025 0.56 0.9675 ;
        RECT 0.435 0.9025 0.5 1.2825 ;
        RECT 0.245 0.265 0.31 0.9675 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 0.56 1.55 ;
        RECT 0.06 1.04 0.125 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.56 0.2 ;
        RECT 0.435 0 0.5 0.415 ;
        RECT 0.06 0 0.125 0.415 ;
    END
  END vss!
END nor2

MACRO oai21
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN oai21 0 0.1 ;
  SIZE 0.75 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.09 0.4975 0.155 0.6325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.395 0.5325 0.46 0.6675 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.595 0.4975 0.66 0.6325 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.245 0.755 0.705 0.82 ;
        RECT 0.435 0.755 0.5 1.2825 ;
        RECT 0.245 0.265 0.31 0.82 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 0.755 1.55 ;
        RECT 0.6275 1.04 0.6925 1.55 ;
        RECT 0.06 1.04 0.125 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.75 0.2 ;
        RECT 0.625 0 0.69 0.415 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.435 0.265 0.5 0.415 ;
      RECT 0.06 0.265 0.125 0.415 ;
    LAYER metal2 ;
      RECT 0.0575 0.47 0.5025 0.54 ;
      RECT 0.4325 0.275 0.5025 0.54 ;
      RECT 0.0575 0.275 0.1275 0.54 ;
    LAYER via1 ;
      RECT 0.435 0.31 0.5 0.375 ;
      RECT 0.06 0.31 0.125 0.375 ;
  END
END oai21

MACRO or2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN or2 0 0.1 ;
  SIZE 0.75 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.57 0.555 0.705 0.62 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2925 0.4975 0.3575 0.6325 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.265 0.125 1.2825 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 0.75 1.55 ;
        RECT 0.25 1.04 0.315 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.75 0.2 ;
        RECT 0.625 0 0.69 0.415 ;
        RECT 0.25 0 0.315 0.415 ;
    END
  END vss!
  OBS
    LAYER metal1 ;
      RECT 0.625 0.875 0.69 1.2825 ;
      RECT 0.2025 0.84 0.2675 0.975 ;
      RECT 0.2025 0.875 0.69 0.94 ;
      RECT 0.435 0.265 0.5 0.94 ;
  END
END or2

MACRO xnor2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN xnor2 0 0.1 ;
  SIZE 1.13 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.625 0.8225 0.8825 0.8875 ;
        RECT 0.8175 0.265 0.8825 0.8875 ;
        RECT 0.625 0.8225 0.69 1.285 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 1.13 1.55 ;
        RECT 1.005 1.0425 1.07 1.55 ;
        RECT 0.435 1.0425 0.5 1.55 ;
        RECT 0.06 1.04 0.125 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 1.13 0.2 ;
        RECT 0.435 0 0.5 0.415 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.0475 0.805 1.0825 0.875 ;
      LAYER metal1 ;
        RECT 0.9475 0.8075 1.0825 0.8725 ;
        RECT 0.0475 0.8075 0.1825 0.8725 ;
      LAYER via1 ;
        RECT 0.0825 0.8075 0.1475 0.8725 ;
        RECT 0.9825 0.8075 1.0475 0.8725 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.3575 0.4975 0.4925 0.5675 ;
      LAYER metal1 ;
        RECT 0.6825 0.5 0.7475 0.635 ;
        RECT 0.3575 0.5 0.7475 0.565 ;
      LAYER via1 ;
        RECT 0.3925 0.5 0.4575 0.565 ;
    END
  END B
  OBS
    LAYER metal1 ;
      RECT 0.2475 0.645 0.3125 1.2825 ;
      RECT 0.48 0.645 0.545 0.78 ;
      RECT 0.06 0.645 0.545 0.71 ;
      RECT 0.06 0.265 0.125 0.71 ;
      RECT 1.005 0.265 1.07 0.415 ;
      RECT 0.6275 0.265 0.6925 0.415 ;
    LAYER metal2 ;
      RECT 1.0025 0.2725 1.0725 0.4075 ;
      RECT 0.625 0.2725 0.695 0.4075 ;
      RECT 0.625 0.2725 1.0725 0.3425 ;
    LAYER via1 ;
      RECT 1.005 0.3075 1.07 0.3725 ;
      RECT 0.6275 0.3075 0.6925 0.3725 ;
  END
END xnor2

MACRO xor2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN xor2 0 0.1 ;
  SIZE 1.13 BY 1.35 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.68 0.6375 0.745 0.7725 ;
        RECT 0.3925 0.6725 0.745 0.7375 ;
        RECT 0.3925 0.6375 0.4575 0.7725 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.8125 0.4725 0.8825 1.2825 ;
        RECT 0.6225 0.4725 0.8825 0.5425 ;
        RECT 0.6225 0.265 0.6925 0.5425 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.35 1.13 1.55 ;
        RECT 0.435 1.0425 0.5 1.55 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 1.13 0.2 ;
        RECT 1.005 0 1.07 0.415 ;
        RECT 0.435 0 0.5 0.415 ;
        RECT 0.06 0 0.125 0.415 ;
    END
  END vss!
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.9725 0.5025 1.0425 0.6375 ;
        RECT 0.0875 0.5375 1.0425 0.6075 ;
        RECT 0.0875 0.5025 0.1575 0.6375 ;
      LAYER metal1 ;
        RECT 0.975 0.5025 1.04 0.6375 ;
        RECT 0.09 0.5025 0.155 0.6375 ;
      LAYER via1 ;
        RECT 0.09 0.5375 0.155 0.6025 ;
        RECT 0.975 0.5375 1.04 0.6025 ;
    END
  END B
  OBS
    LAYER metal1 ;
      RECT 0.06 0.9075 0.125 1.2825 ;
      RECT 0.06 0.9075 0.5825 0.9725 ;
      RECT 0.245 0.265 0.31 0.9725 ;
      RECT 1.005 1.0425 1.07 1.2825 ;
      RECT 0.625 1.0425 0.69 1.2825 ;
    LAYER metal2 ;
      RECT 1.0025 0.9525 1.0725 1.23 ;
      RECT 0.6225 0.9525 0.6925 1.23 ;
      RECT 0.6225 0.9525 1.0725 1.0225 ;
    LAYER via1 ;
      RECT 1.005 1.13 1.07 1.195 ;
      RECT 0.625 1.13 0.69 1.195 ;
  END
END xor2

END LIBRARY
